//////////////////////////////////////////////////////////////////////
// Created by SmartDesign Tue Mar 29 05:35:45 2022
// Version: v2021.2 2021.2.0.11
//////////////////////////////////////////////////////////////////////

`timescale 1ns / 100ps

//////////////////////////////////////////////////////////////////////
// Component Description (Tcl) 
//////////////////////////////////////////////////////////////////////
/*
# Exporting Component Description of PF_DDR4_SS_DDRPHY_BLK to TCL
# Family: PolarFire
# Part Number: MPF100T-1FCVG484I
# Create and Configure the core component PF_DDR4_SS_DDRPHY_BLK
create_and_configure_core -core_vlnv {Actel:SystemBuilder:PF_DDR4PHY:2.4.104} -component_name {PF_DDR4_SS_DDRPHY_BLK} -params {\
"IOG_CLOCK_RATIO:4" \
"IOG_NUM_BCLKS:1" \
"IOG_WRITE_LEVELING:1" \
"PIPELINE:true" \
"SDRAM_BG_ADDR_WIDTH:2" \
"SDRAM_DATA_RATE:1600.0" \
"SDRAM_DATA_WIDTH:32" \
"SDRAM_DM_MODE:1" \
"SDRAM_NB_RANKS:1" \
"SDRAM_NUM_CLK_OUTS:1" \
"SDRAM_PARITY_ALERT:0" \
"SDRAM_ROW_ADDR_WIDTH:15" \
"SDRAM_TYPE:0" \
"SHIELD_ENABLED:true" \
"SIMULATION_MODE:FAST" }
# Exporting Component Description of PF_DDR4_SS_DDRPHY_BLK to TCL done
*/

// PF_DDR4_SS_DDRPHY_BLK
module PF_DDR4_SS_DDRPHY_BLK(
    // Inputs
    ADDR_VCOPHS_OFFSET,
    ADDR_WAIT_COUNT,
    BCLK_VCOPHS_OFFSET,
    CAL_INIT_ACK,
    CAL_L_BUSY,
    CAL_L_DATAOUT,
    CAL_L_D_REQ,
    CAL_L_R_VALID,
    CTRLR_READY_IN,
    DFI_ACT_N_P0,
    DFI_ACT_N_P1,
    DFI_ACT_N_P2,
    DFI_ACT_N_P3,
    DFI_ADDRESS_P0,
    DFI_ADDRESS_P1,
    DFI_ADDRESS_P2,
    DFI_ADDRESS_P3,
    DFI_BANK_P0,
    DFI_BANK_P1,
    DFI_BANK_P2,
    DFI_BANK_P3,
    DFI_BG_P0,
    DFI_BG_P1,
    DFI_BG_P2,
    DFI_BG_P3,
    DFI_CALVL_BG_PATTERN,
    DFI_CALVL_CAPTURE,
    DFI_CALVL_EN,
    DFI_CALVL_START,
    DFI_CALVL_TRN_COMMAND,
    DFI_CAS_N_P0,
    DFI_CAS_N_P1,
    DFI_CAS_N_P2,
    DFI_CAS_N_P3,
    DFI_CKE_P0,
    DFI_CKE_P1,
    DFI_CKE_P2,
    DFI_CKE_P3,
    DFI_CS_N_P0,
    DFI_CS_N_P1,
    DFI_CS_N_P2,
    DFI_CS_N_P3,
    DFI_CTRLR_BUSY,
    DFI_CTRLUPD_REQ,
    DFI_INIT_START,
    DFI_LVL_PATTERN,
    DFI_LVL_PERIODIC,
    DFI_ODT_P0,
    DFI_ODT_P1,
    DFI_ODT_P2,
    DFI_ODT_P3,
    DFI_PHYUPD_ACK,
    DFI_RAS_N_P0,
    DFI_RAS_N_P1,
    DFI_RAS_N_P2,
    DFI_RAS_N_P3,
    DFI_RDDATA_CS_N_P0,
    DFI_RDDATA_CS_N_P1,
    DFI_RDDATA_CS_N_P2,
    DFI_RDDATA_CS_N_P3,
    DFI_RDDATA_EN_P0,
    DFI_RDDATA_EN_P1,
    DFI_RDDATA_EN_P2,
    DFI_RDDATA_EN_P3,
    DFI_RDLVL_CS_N,
    DFI_RDLVL_EN,
    DFI_RDLVL_GATE_EN,
    DFI_RESET_N_P0,
    DFI_RESET_N_P1,
    DFI_RESET_N_P2,
    DFI_RESET_N_P3,
    DFI_WE_N_P0,
    DFI_WE_N_P1,
    DFI_WE_N_P2,
    DFI_WE_N_P3,
    DFI_WRDATA_CS_N_P0,
    DFI_WRDATA_CS_N_P1,
    DFI_WRDATA_CS_N_P2,
    DFI_WRDATA_CS_N_P3,
    DFI_WRDATA_EN_P0,
    DFI_WRDATA_EN_P1,
    DFI_WRDATA_EN_P2,
    DFI_WRDATA_EN_P3,
    DFI_WRDATA_MASK_P0,
    DFI_WRDATA_MASK_P1,
    DFI_WRDATA_MASK_P2,
    DFI_WRDATA_MASK_P3,
    DFI_WRDATA_P0,
    DFI_WRDATA_P1,
    DFI_WRDATA_P2,
    DFI_WRDATA_P3,
    DFI_WRLVL_CS_N,
    DFI_WRLVL_EN,
    DFI_WRLVL_STROBE,
    DLL_CODE,
    DLL_DLY_DIFF,
    HS_IO_CLK,
    HS_IO_CLK_270,
    PADDR,
    PCLK,
    PENABLE,
    PLL_LOCK,
    PSEL,
    PWDATA,
    PWRITE,
    RDGATE_MIN_READS_THRESHOLD,
    REF_CLK,
    SKIP_BCLK_TRN,
    SKIP_CA_TRN,
    SKIP_DQSW_TRN,
    SKIP_RDLVL_TRN,
    SKIP_VREF_TRAINING,
    SKIP_WRLVL_TRN,
    SYS_CLK,
    SYS_RST_N,
    VREF_MR6_VALUE,
    WRCAL_WRITE_COUNTER_VALUE,
    WRLVL_TAP_OFFSET,
    // Outputs
    A,
    ACT_N,
    BA,
    BG,
    CAL_INIT_CS,
    CAL_INIT_MR_ADDR,
    CAL_INIT_MR_WR_DATA,
    CAL_INIT_MR_WR_MASK,
    CAL_INIT_MR_W_REQ,
    CAL_L_DATAIN,
    CAL_L_DM_IN,
    CAL_L_R_REQ,
    CAL_L_W_REQ,
    CAL_SELECT,
    CAS_N,
    CK0,
    CK0_N,
    CKE,
    CODE_UPDATE,
    CS_N,
    CTRLR_READY_OUT,
    DFI_CALVL_RESP,
    DFI_CALVL_TRAIN_DONE,
    DFI_CTRLUPD_ACK,
    DFI_INIT_COMPLETE,
    DFI_PHYUPD_REQ,
    DFI_PHYUPD_TYPE,
    DFI_RDDATA_VALID_W0,
    DFI_RDDATA_VALID_W1,
    DFI_RDDATA_VALID_W2,
    DFI_RDDATA_VALID_W3,
    DFI_RDDATA_W0,
    DFI_RDDATA_W1,
    DFI_RDDATA_W2,
    DFI_RDDATA_W3,
    DFI_RDLVL_RESP,
    DFI_TRAINING_COMPLETE,
    DFI_WRLVL_RESP,
    DM_N,
    ITER_COUNT,
    LOADPHS_B,
    ODT,
    PRDATA,
    PREADY,
    RAS_N,
    RESET_N,
    SHIELD0,
    SHIELD1,
    SHIELD2,
    SHIELD3,
    SYNC_SYS_RST_N,
    VCO_PHSEL_BCLK90_SEL,
    VCO_PHSEL_BCLK_SEL,
    VCO_PHSEL_REFCLK_SEL,
    VCO_PHSEL_ROTATE,
    WE_N,
    // Inouts
    DQ,
    DQS,
    DQS_N
);

//--------------------------------------------------------------------
// Input
//--------------------------------------------------------------------
input  [2:0]   ADDR_VCOPHS_OFFSET;
input  [9:0]   ADDR_WAIT_COUNT;
input  [2:0]   BCLK_VCOPHS_OFFSET;
input          CAL_INIT_ACK;
input          CAL_L_BUSY;
input  [255:0] CAL_L_DATAOUT;
input          CAL_L_D_REQ;
input          CAL_L_R_VALID;
input          CTRLR_READY_IN;
input          DFI_ACT_N_P0;
input          DFI_ACT_N_P1;
input          DFI_ACT_N_P2;
input          DFI_ACT_N_P3;
input  [16:0]  DFI_ADDRESS_P0;
input  [16:0]  DFI_ADDRESS_P1;
input  [16:0]  DFI_ADDRESS_P2;
input  [16:0]  DFI_ADDRESS_P3;
input  [1:0]   DFI_BANK_P0;
input  [1:0]   DFI_BANK_P1;
input  [1:0]   DFI_BANK_P2;
input  [1:0]   DFI_BANK_P3;
input  [1:0]   DFI_BG_P0;
input  [1:0]   DFI_BG_P1;
input  [1:0]   DFI_BG_P2;
input  [1:0]   DFI_BG_P3;
input  [19:0]  DFI_CALVL_BG_PATTERN;
input          DFI_CALVL_CAPTURE;
input          DFI_CALVL_EN;
input          DFI_CALVL_START;
input  [19:0]  DFI_CALVL_TRN_COMMAND;
input          DFI_CAS_N_P0;
input          DFI_CAS_N_P1;
input          DFI_CAS_N_P2;
input          DFI_CAS_N_P3;
input  [0:0]   DFI_CKE_P0;
input  [0:0]   DFI_CKE_P1;
input  [0:0]   DFI_CKE_P2;
input  [0:0]   DFI_CKE_P3;
input  [0:0]   DFI_CS_N_P0;
input  [0:0]   DFI_CS_N_P1;
input  [0:0]   DFI_CS_N_P2;
input  [0:0]   DFI_CS_N_P3;
input          DFI_CTRLR_BUSY;
input          DFI_CTRLUPD_REQ;
input          DFI_INIT_START;
input  [3:0]   DFI_LVL_PATTERN;
input          DFI_LVL_PERIODIC;
input  [0:0]   DFI_ODT_P0;
input  [0:0]   DFI_ODT_P1;
input  [0:0]   DFI_ODT_P2;
input  [0:0]   DFI_ODT_P3;
input          DFI_PHYUPD_ACK;
input          DFI_RAS_N_P0;
input          DFI_RAS_N_P1;
input          DFI_RAS_N_P2;
input          DFI_RAS_N_P3;
input  [0:0]   DFI_RDDATA_CS_N_P0;
input  [0:0]   DFI_RDDATA_CS_N_P1;
input  [0:0]   DFI_RDDATA_CS_N_P2;
input  [0:0]   DFI_RDDATA_CS_N_P3;
input  [31:0]  DFI_RDDATA_EN_P0;
input  [31:0]  DFI_RDDATA_EN_P1;
input  [31:0]  DFI_RDDATA_EN_P2;
input  [31:0]  DFI_RDDATA_EN_P3;
input  [0:0]   DFI_RDLVL_CS_N;
input          DFI_RDLVL_EN;
input          DFI_RDLVL_GATE_EN;
input          DFI_RESET_N_P0;
input          DFI_RESET_N_P1;
input          DFI_RESET_N_P2;
input          DFI_RESET_N_P3;
input          DFI_WE_N_P0;
input          DFI_WE_N_P1;
input          DFI_WE_N_P2;
input          DFI_WE_N_P3;
input  [0:0]   DFI_WRDATA_CS_N_P0;
input  [0:0]   DFI_WRDATA_CS_N_P1;
input  [0:0]   DFI_WRDATA_CS_N_P2;
input  [0:0]   DFI_WRDATA_CS_N_P3;
input  [31:0]  DFI_WRDATA_EN_P0;
input  [31:0]  DFI_WRDATA_EN_P1;
input  [31:0]  DFI_WRDATA_EN_P2;
input  [31:0]  DFI_WRDATA_EN_P3;
input  [7:0]   DFI_WRDATA_MASK_P0;
input  [7:0]   DFI_WRDATA_MASK_P1;
input  [7:0]   DFI_WRDATA_MASK_P2;
input  [7:0]   DFI_WRDATA_MASK_P3;
input  [63:0]  DFI_WRDATA_P0;
input  [63:0]  DFI_WRDATA_P1;
input  [63:0]  DFI_WRDATA_P2;
input  [63:0]  DFI_WRDATA_P3;
input  [0:0]   DFI_WRLVL_CS_N;
input          DFI_WRLVL_EN;
input          DFI_WRLVL_STROBE;
input  [7:0]   DLL_CODE;
input          DLL_DLY_DIFF;
input          HS_IO_CLK;
input          HS_IO_CLK_270;
input  [15:0]  PADDR;
input          PCLK;
input          PENABLE;
input          PLL_LOCK;
input          PSEL;
input  [7:0]   PWDATA;
input          PWRITE;
input  [9:0]   RDGATE_MIN_READS_THRESHOLD;
input          REF_CLK;
input          SKIP_BCLK_TRN;
input          SKIP_CA_TRN;
input          SKIP_DQSW_TRN;
input          SKIP_RDLVL_TRN;
input          SKIP_VREF_TRAINING;
input          SKIP_WRLVL_TRN;
input          SYS_CLK;
input          SYS_RST_N;
input  [6:0]   VREF_MR6_VALUE;
input  [7:0]   WRCAL_WRITE_COUNTER_VALUE;
input  [6:0]   WRLVL_TAP_OFFSET;
//--------------------------------------------------------------------
// Output
//--------------------------------------------------------------------
output [13:0]  A;
output         ACT_N;
output [1:0]   BA;
output [1:0]   BG;
output [1:0]   CAL_INIT_CS;
output [7:0]   CAL_INIT_MR_ADDR;
output [17:0]  CAL_INIT_MR_WR_DATA;
output [17:0]  CAL_INIT_MR_WR_MASK;
output         CAL_INIT_MR_W_REQ;
output [255:0] CAL_L_DATAIN;
output [31:0]  CAL_L_DM_IN;
output         CAL_L_R_REQ;
output         CAL_L_W_REQ;
output         CAL_SELECT;
output         CAS_N;
output         CK0;
output         CK0_N;
output         CKE;
output         CODE_UPDATE;
output         CS_N;
output         CTRLR_READY_OUT;
output [1:0]   DFI_CALVL_RESP;
output         DFI_CALVL_TRAIN_DONE;
output         DFI_CTRLUPD_ACK;
output         DFI_INIT_COMPLETE;
output         DFI_PHYUPD_REQ;
output [1:0]   DFI_PHYUPD_TYPE;
output [3:0]   DFI_RDDATA_VALID_W0;
output [3:0]   DFI_RDDATA_VALID_W1;
output [3:0]   DFI_RDDATA_VALID_W2;
output [3:0]   DFI_RDDATA_VALID_W3;
output [63:0]  DFI_RDDATA_W0;
output [63:0]  DFI_RDDATA_W1;
output [63:0]  DFI_RDDATA_W2;
output [63:0]  DFI_RDDATA_W3;
output [3:0]   DFI_RDLVL_RESP;
output         DFI_TRAINING_COMPLETE;
output [3:0]   DFI_WRLVL_RESP;
output [3:0]   DM_N;
output [3:0]   ITER_COUNT;
output [0:0]   LOADPHS_B;
output         ODT;
output [7:0]   PRDATA;
output         PREADY;
output         RAS_N;
output         RESET_N;
output         SHIELD0;
output         SHIELD1;
output         SHIELD2;
output         SHIELD3;
output         SYNC_SYS_RST_N;
output [0:0]   VCO_PHSEL_BCLK90_SEL;
output [0:0]   VCO_PHSEL_BCLK_SEL;
output         VCO_PHSEL_REFCLK_SEL;
output [0:0]   VCO_PHSEL_ROTATE;
output         WE_N;
//--------------------------------------------------------------------
// Inout
//--------------------------------------------------------------------
inout  [31:0]  DQ;
inout  [3:0]   DQS;
inout  [3:0]   DQS_N;
//--------------------------------------------------------------------
// Nets
//--------------------------------------------------------------------
wire   [0:0]     A_net_0;
wire   [1:1]     A_0;
wire   [2:2]     A_1;
wire   [3:3]     A_2;
wire   [4:4]     A_3;
wire   [5:5]     A_4;
wire   [6:6]     A_5;
wire   [7:7]     A_6;
wire   [8:8]     A_7;
wire   [9:9]     A_8;
wire   [10:10]   A_9;
wire   [11:11]   A_10;
wire             A_11;
wire   [0:0]     A_12;
wire   [0:0]     ACT_N_net_0;
wire   [2:0]     ADDR_VCOPHS_OFFSET;
wire   [9:0]     ADDR_WAIT_COUNT;
wire   [15:0]    PADDR;
wire             PENABLE;
wire   [7:0]     APB_DEBUG_PRDATA;
wire             APB_DEBUG_PREADY;
wire             PSEL;
wire   [7:0]     PWDATA;
wire             PWRITE;
wire   [1:0]     BA_net_0;
wire   [2:0]     BCLK_VCOPHS_OFFSET;
wire   [1:0]     BG_net_0;
wire             CAL_INIT_ACK;
wire   [1:0]     CAL_INIT_CS_net_0;
wire   [7:0]     CAL_INIT_MR_ADDR_net_0;
wire             CAL_INIT_MR_W_REQ_net_0;
wire   [17:0]    CAL_INIT_MR_WR_DATA_net_0;
wire   [17:0]    CAL_INIT_MR_WR_MASK_net_0;
wire             CAL_L_BUSY;
wire             CAL_L_D_REQ;
wire   [255:0]   CAL_L_DATAIN_net_0;
wire   [255:0]   CAL_L_DATAOUT;
wire   [31:0]    CAL_L_DM_IN_net_0;
wire             CAL_L_R_REQ_net_0;
wire             CAL_L_R_VALID;
wire             CAL_L_W_REQ_net_0;
wire             CAL_SELECT_net_0;
wire   [0:0]     CAS_N_net_0;
wire             CK0_net_0;
wire             CK0_N_net_0;
wire   [0:0]     CKE_net_0;
wire             CLKINT_CMD_Y;
wire             CODE_UPDATE_net_0;
wire   [0:0]     CS_N_net_0;
wire             CTRLR_READY_IN;
wire             CTRLR_READY_OUT_net_0;
wire             DFI_ACT_N_P0;
wire             DFI_ACT_N_P1;
wire             DFI_ACT_N_P2;
wire             DFI_ACT_N_P3;
wire   [0:0]     DFI_ADDRESS_P0_slice_0;
wire   [1:1]     DFI_ADDRESS_P0_slice_1;
wire   [2:2]     DFI_ADDRESS_P0_slice_2;
wire   [3:3]     DFI_ADDRESS_P0_slice_3;
wire   [4:4]     DFI_ADDRESS_P0_slice_4;
wire   [5:5]     DFI_ADDRESS_P0_slice_5;
wire   [6:6]     DFI_ADDRESS_P0_slice_6;
wire   [7:7]     DFI_ADDRESS_P0_slice_7;
wire   [8:8]     DFI_ADDRESS_P0_slice_8;
wire   [9:9]     DFI_ADDRESS_P0_slice_9;
wire   [10:10]   DFI_ADDRESS_P0_slice_10;
wire   [11:11]   DFI_ADDRESS_P0_slice_11;
wire   [12:12]   DFI_ADDRESS_P0_slice_12;
wire   [13:13]   DFI_ADDRESS_P0_slice_13;
wire   [0:0]     DFI_ADDRESS_P1_slice_0;
wire   [1:1]     DFI_ADDRESS_P1_slice_1;
wire   [2:2]     DFI_ADDRESS_P1_slice_2;
wire   [3:3]     DFI_ADDRESS_P1_slice_3;
wire   [4:4]     DFI_ADDRESS_P1_slice_4;
wire   [5:5]     DFI_ADDRESS_P1_slice_5;
wire   [6:6]     DFI_ADDRESS_P1_slice_6;
wire   [7:7]     DFI_ADDRESS_P1_slice_7;
wire   [8:8]     DFI_ADDRESS_P1_slice_8;
wire   [9:9]     DFI_ADDRESS_P1_slice_9;
wire   [10:10]   DFI_ADDRESS_P1_slice_10;
wire   [11:11]   DFI_ADDRESS_P1_slice_11;
wire   [12:12]   DFI_ADDRESS_P1_slice_12;
wire   [13:13]   DFI_ADDRESS_P1_slice_13;
wire   [0:0]     DFI_ADDRESS_P2_slice_0;
wire   [1:1]     DFI_ADDRESS_P2_slice_1;
wire   [2:2]     DFI_ADDRESS_P2_slice_2;
wire   [3:3]     DFI_ADDRESS_P2_slice_3;
wire   [4:4]     DFI_ADDRESS_P2_slice_4;
wire   [5:5]     DFI_ADDRESS_P2_slice_5;
wire   [6:6]     DFI_ADDRESS_P2_slice_6;
wire   [7:7]     DFI_ADDRESS_P2_slice_7;
wire   [8:8]     DFI_ADDRESS_P2_slice_8;
wire   [9:9]     DFI_ADDRESS_P2_slice_9;
wire   [10:10]   DFI_ADDRESS_P2_slice_10;
wire   [11:11]   DFI_ADDRESS_P2_slice_11;
wire   [12:12]   DFI_ADDRESS_P2_slice_12;
wire   [13:13]   DFI_ADDRESS_P2_slice_13;
wire   [0:0]     DFI_ADDRESS_P3_slice_0;
wire   [1:1]     DFI_ADDRESS_P3_slice_1;
wire   [2:2]     DFI_ADDRESS_P3_slice_2;
wire   [3:3]     DFI_ADDRESS_P3_slice_3;
wire   [4:4]     DFI_ADDRESS_P3_slice_4;
wire   [5:5]     DFI_ADDRESS_P3_slice_5;
wire   [6:6]     DFI_ADDRESS_P3_slice_6;
wire   [7:7]     DFI_ADDRESS_P3_slice_7;
wire   [8:8]     DFI_ADDRESS_P3_slice_8;
wire   [9:9]     DFI_ADDRESS_P3_slice_9;
wire   [10:10]   DFI_ADDRESS_P3_slice_10;
wire   [11:11]   DFI_ADDRESS_P3_slice_11;
wire   [12:12]   DFI_ADDRESS_P3_slice_12;
wire   [13:13]   DFI_ADDRESS_P3_slice_13;
wire   [0:0]     DFI_BANK_P0_slice_0;
wire   [1:1]     DFI_BANK_P0_slice_1;
wire   [0:0]     DFI_BANK_P1_slice_0;
wire   [1:1]     DFI_BANK_P1_slice_1;
wire   [0:0]     DFI_BANK_P2_slice_0;
wire   [1:1]     DFI_BANK_P2_slice_1;
wire   [0:0]     DFI_BANK_P3_slice_0;
wire   [1:1]     DFI_BANK_P3_slice_1;
wire   [0:0]     DFI_BG_P0_slice_0;
wire   [1:1]     DFI_BG_P0_slice_1;
wire   [0:0]     DFI_BG_P1_slice_0;
wire   [1:1]     DFI_BG_P1_slice_1;
wire   [0:0]     DFI_BG_P2_slice_0;
wire   [1:1]     DFI_BG_P2_slice_1;
wire   [0:0]     DFI_BG_P3_slice_0;
wire   [1:1]     DFI_BG_P3_slice_1;
wire             DFI_CAS_N_P0;
wire             DFI_CAS_N_P1;
wire             DFI_CAS_N_P2;
wire             DFI_CAS_N_P3;
wire   [0:0]     DFI_CKE_P0;
wire   [0:0]     DFI_CKE_P1;
wire   [0:0]     DFI_CKE_P2;
wire   [0:0]     DFI_CKE_P3;
wire   [0:0]     DFI_CS_N_P0;
wire   [0:0]     DFI_CS_N_P1;
wire   [0:0]     DFI_CS_N_P2;
wire   [0:0]     DFI_CS_N_P3;
wire             DFI_CTRLUPD_REQ;
wire             DFI_INIT_COMPLETE_net_0;
wire             DFI_INIT_START;
wire   [0:0]     DFI_ODT_P0;
wire   [0:0]     DFI_ODT_P1;
wire   [0:0]     DFI_ODT_P2;
wire   [0:0]     DFI_ODT_P3;
wire             DFI_RAS_N_P0;
wire             DFI_RAS_N_P1;
wire             DFI_RAS_N_P2;
wire             DFI_RAS_N_P3;
wire   [0:0]     DFI_RDDATA_CS_N_P0;
wire   [0:0]     DFI_RDDATA_CS_N_P1;
wire   [0:0]     DFI_RDDATA_CS_N_P2;
wire   [0:0]     DFI_RDDATA_CS_N_P3;
wire   [0:0]     DFI_RDDATA_EN_P0_slice_0;
wire   [0:0]     DFI_RDDATA_EN_P1_slice_0;
wire   [0:0]     DFI_RDDATA_EN_P2_slice_0;
wire   [0:0]     DFI_RDDATA_EN_P3_slice_0;
wire             DFI_RDDATA_VALID_W0_net_0;
wire             DFI_RDDATA_VALID_W1_net_0;
wire             DFI_RDDATA_VALID_W2_net_0;
wire             DFI_RDDATA_VALID_W3_net_0;
wire   [63:0]    DFI_RDDATA_W0_net_0;
wire   [63:0]    DFI_RDDATA_W1_net_0;
wire   [63:0]    DFI_RDDATA_W2_net_0;
wire   [63:0]    DFI_RDDATA_W3_net_0;
wire   [0:0]     DFI_RDLVL_CS_N;
wire             DFI_RDLVL_EN;
wire             DFI_RDLVL_GATE_EN;
wire   [3:0]     DFI_RDLVL_RESP_net_0;
wire             DFI_RESET_N_P0;
wire             DFI_RESET_N_P1;
wire             DFI_RESET_N_P2;
wire             DFI_RESET_N_P3;
wire             DFI_TRAINING_COMPLETE_net_0;
wire             DFI_WE_N_P0;
wire             DFI_WE_N_P1;
wire             DFI_WE_N_P2;
wire             DFI_WE_N_P3;
wire   [0:0]     DFI_WRDATA_CS_N_P0;
wire   [0:0]     DFI_WRDATA_CS_N_P1;
wire   [0:0]     DFI_WRDATA_CS_N_P2;
wire   [0:0]     DFI_WRDATA_CS_N_P3;
wire   [0:0]     DFI_WRDATA_EN_P0_slice_0;
wire   [0:0]     DFI_WRDATA_EN_P1_slice_0;
wire   [0:0]     DFI_WRDATA_EN_P2_slice_0;
wire   [0:0]     DFI_WRDATA_EN_P3_slice_0;
wire   [0:0]     DFI_WRDATA_MASK_P0_slice_0;
wire   [4:4]     DFI_WRDATA_MASK_P0_slice_1;
wire   [1:1]     DFI_WRDATA_MASK_P0_slice_2;
wire   [5:5]     DFI_WRDATA_MASK_P0_slice_3;
wire   [2:2]     DFI_WRDATA_MASK_P0_slice_4;
wire   [6:6]     DFI_WRDATA_MASK_P0_slice_5;
wire   [3:3]     DFI_WRDATA_MASK_P0_slice_6;
wire   [7:7]     DFI_WRDATA_MASK_P0_slice_7;
wire   [0:0]     DFI_WRDATA_MASK_P1_slice_0;
wire   [4:4]     DFI_WRDATA_MASK_P1_slice_1;
wire   [1:1]     DFI_WRDATA_MASK_P1_slice_2;
wire   [5:5]     DFI_WRDATA_MASK_P1_slice_3;
wire   [2:2]     DFI_WRDATA_MASK_P1_slice_4;
wire   [6:6]     DFI_WRDATA_MASK_P1_slice_5;
wire   [3:3]     DFI_WRDATA_MASK_P1_slice_6;
wire   [7:7]     DFI_WRDATA_MASK_P1_slice_7;
wire   [0:0]     DFI_WRDATA_MASK_P2_slice_0;
wire   [4:4]     DFI_WRDATA_MASK_P2_slice_1;
wire   [1:1]     DFI_WRDATA_MASK_P2_slice_2;
wire   [5:5]     DFI_WRDATA_MASK_P2_slice_3;
wire   [2:2]     DFI_WRDATA_MASK_P2_slice_4;
wire   [6:6]     DFI_WRDATA_MASK_P2_slice_5;
wire   [3:3]     DFI_WRDATA_MASK_P2_slice_6;
wire   [7:7]     DFI_WRDATA_MASK_P2_slice_7;
wire   [0:0]     DFI_WRDATA_MASK_P3_slice_0;
wire   [4:4]     DFI_WRDATA_MASK_P3_slice_1;
wire   [1:1]     DFI_WRDATA_MASK_P3_slice_2;
wire   [5:5]     DFI_WRDATA_MASK_P3_slice_3;
wire   [2:2]     DFI_WRDATA_MASK_P3_slice_4;
wire   [6:6]     DFI_WRDATA_MASK_P3_slice_5;
wire   [3:3]     DFI_WRDATA_MASK_P3_slice_6;
wire   [7:7]     DFI_WRDATA_MASK_P3_slice_7;
wire   [0:0]     DFI_WRDATA_P0_slice_0;
wire   [32:32]   DFI_WRDATA_P0_slice_1;
wire   [1:1]     DFI_WRDATA_P0_slice_2;
wire   [33:33]   DFI_WRDATA_P0_slice_3;
wire   [2:2]     DFI_WRDATA_P0_slice_4;
wire   [34:34]   DFI_WRDATA_P0_slice_5;
wire   [3:3]     DFI_WRDATA_P0_slice_6;
wire   [35:35]   DFI_WRDATA_P0_slice_7;
wire   [4:4]     DFI_WRDATA_P0_slice_8;
wire   [36:36]   DFI_WRDATA_P0_slice_9;
wire   [5:5]     DFI_WRDATA_P0_slice_10;
wire   [37:37]   DFI_WRDATA_P0_slice_11;
wire   [6:6]     DFI_WRDATA_P0_slice_12;
wire   [38:38]   DFI_WRDATA_P0_slice_13;
wire   [7:7]     DFI_WRDATA_P0_slice_14;
wire   [39:39]   DFI_WRDATA_P0_slice_15;
wire   [8:8]     DFI_WRDATA_P0_slice_16;
wire   [40:40]   DFI_WRDATA_P0_slice_17;
wire   [9:9]     DFI_WRDATA_P0_slice_18;
wire   [41:41]   DFI_WRDATA_P0_slice_19;
wire   [10:10]   DFI_WRDATA_P0_slice_20;
wire   [42:42]   DFI_WRDATA_P0_slice_21;
wire   [11:11]   DFI_WRDATA_P0_slice_22;
wire   [43:43]   DFI_WRDATA_P0_slice_23;
wire   [12:12]   DFI_WRDATA_P0_slice_24;
wire   [44:44]   DFI_WRDATA_P0_slice_25;
wire   [13:13]   DFI_WRDATA_P0_slice_26;
wire   [45:45]   DFI_WRDATA_P0_slice_27;
wire   [14:14]   DFI_WRDATA_P0_slice_28;
wire   [46:46]   DFI_WRDATA_P0_slice_29;
wire   [15:15]   DFI_WRDATA_P0_slice_30;
wire   [47:47]   DFI_WRDATA_P0_slice_31;
wire   [16:16]   DFI_WRDATA_P0_slice_32;
wire   [48:48]   DFI_WRDATA_P0_slice_33;
wire   [17:17]   DFI_WRDATA_P0_slice_34;
wire   [49:49]   DFI_WRDATA_P0_slice_35;
wire   [18:18]   DFI_WRDATA_P0_slice_36;
wire   [50:50]   DFI_WRDATA_P0_slice_37;
wire   [19:19]   DFI_WRDATA_P0_slice_38;
wire   [51:51]   DFI_WRDATA_P0_slice_39;
wire   [20:20]   DFI_WRDATA_P0_slice_40;
wire   [52:52]   DFI_WRDATA_P0_slice_41;
wire   [21:21]   DFI_WRDATA_P0_slice_42;
wire   [53:53]   DFI_WRDATA_P0_slice_43;
wire   [22:22]   DFI_WRDATA_P0_slice_44;
wire   [54:54]   DFI_WRDATA_P0_slice_45;
wire   [23:23]   DFI_WRDATA_P0_slice_46;
wire   [55:55]   DFI_WRDATA_P0_slice_47;
wire   [24:24]   DFI_WRDATA_P0_slice_48;
wire   [56:56]   DFI_WRDATA_P0_slice_49;
wire   [25:25]   DFI_WRDATA_P0_slice_50;
wire   [57:57]   DFI_WRDATA_P0_slice_51;
wire   [26:26]   DFI_WRDATA_P0_slice_52;
wire   [58:58]   DFI_WRDATA_P0_slice_53;
wire   [27:27]   DFI_WRDATA_P0_slice_54;
wire   [59:59]   DFI_WRDATA_P0_slice_55;
wire   [28:28]   DFI_WRDATA_P0_slice_56;
wire   [60:60]   DFI_WRDATA_P0_slice_57;
wire   [29:29]   DFI_WRDATA_P0_slice_58;
wire   [61:61]   DFI_WRDATA_P0_slice_59;
wire   [30:30]   DFI_WRDATA_P0_slice_60;
wire   [62:62]   DFI_WRDATA_P0_slice_61;
wire   [31:31]   DFI_WRDATA_P0_slice_62;
wire   [63:63]   DFI_WRDATA_P0_slice_63;
wire   [0:0]     DFI_WRDATA_P1_slice_0;
wire   [32:32]   DFI_WRDATA_P1_slice_1;
wire   [1:1]     DFI_WRDATA_P1_slice_2;
wire   [33:33]   DFI_WRDATA_P1_slice_3;
wire   [2:2]     DFI_WRDATA_P1_slice_4;
wire   [34:34]   DFI_WRDATA_P1_slice_5;
wire   [3:3]     DFI_WRDATA_P1_slice_6;
wire   [35:35]   DFI_WRDATA_P1_slice_7;
wire   [4:4]     DFI_WRDATA_P1_slice_8;
wire   [36:36]   DFI_WRDATA_P1_slice_9;
wire   [5:5]     DFI_WRDATA_P1_slice_10;
wire   [37:37]   DFI_WRDATA_P1_slice_11;
wire   [6:6]     DFI_WRDATA_P1_slice_12;
wire   [38:38]   DFI_WRDATA_P1_slice_13;
wire   [7:7]     DFI_WRDATA_P1_slice_14;
wire   [39:39]   DFI_WRDATA_P1_slice_15;
wire   [8:8]     DFI_WRDATA_P1_slice_16;
wire   [40:40]   DFI_WRDATA_P1_slice_17;
wire   [9:9]     DFI_WRDATA_P1_slice_18;
wire   [41:41]   DFI_WRDATA_P1_slice_19;
wire   [10:10]   DFI_WRDATA_P1_slice_20;
wire   [42:42]   DFI_WRDATA_P1_slice_21;
wire   [11:11]   DFI_WRDATA_P1_slice_22;
wire   [43:43]   DFI_WRDATA_P1_slice_23;
wire   [12:12]   DFI_WRDATA_P1_slice_24;
wire   [44:44]   DFI_WRDATA_P1_slice_25;
wire   [13:13]   DFI_WRDATA_P1_slice_26;
wire   [45:45]   DFI_WRDATA_P1_slice_27;
wire   [14:14]   DFI_WRDATA_P1_slice_28;
wire   [46:46]   DFI_WRDATA_P1_slice_29;
wire   [15:15]   DFI_WRDATA_P1_slice_30;
wire   [47:47]   DFI_WRDATA_P1_slice_31;
wire   [16:16]   DFI_WRDATA_P1_slice_32;
wire   [48:48]   DFI_WRDATA_P1_slice_33;
wire   [17:17]   DFI_WRDATA_P1_slice_34;
wire   [49:49]   DFI_WRDATA_P1_slice_35;
wire   [18:18]   DFI_WRDATA_P1_slice_36;
wire   [50:50]   DFI_WRDATA_P1_slice_37;
wire   [19:19]   DFI_WRDATA_P1_slice_38;
wire   [51:51]   DFI_WRDATA_P1_slice_39;
wire   [20:20]   DFI_WRDATA_P1_slice_40;
wire   [52:52]   DFI_WRDATA_P1_slice_41;
wire   [21:21]   DFI_WRDATA_P1_slice_42;
wire   [53:53]   DFI_WRDATA_P1_slice_43;
wire   [22:22]   DFI_WRDATA_P1_slice_44;
wire   [54:54]   DFI_WRDATA_P1_slice_45;
wire   [23:23]   DFI_WRDATA_P1_slice_46;
wire   [55:55]   DFI_WRDATA_P1_slice_47;
wire   [24:24]   DFI_WRDATA_P1_slice_48;
wire   [56:56]   DFI_WRDATA_P1_slice_49;
wire   [25:25]   DFI_WRDATA_P1_slice_50;
wire   [57:57]   DFI_WRDATA_P1_slice_51;
wire   [26:26]   DFI_WRDATA_P1_slice_52;
wire   [58:58]   DFI_WRDATA_P1_slice_53;
wire   [27:27]   DFI_WRDATA_P1_slice_54;
wire   [59:59]   DFI_WRDATA_P1_slice_55;
wire   [28:28]   DFI_WRDATA_P1_slice_56;
wire   [60:60]   DFI_WRDATA_P1_slice_57;
wire   [29:29]   DFI_WRDATA_P1_slice_58;
wire   [61:61]   DFI_WRDATA_P1_slice_59;
wire   [30:30]   DFI_WRDATA_P1_slice_60;
wire   [62:62]   DFI_WRDATA_P1_slice_61;
wire   [31:31]   DFI_WRDATA_P1_slice_62;
wire   [63:63]   DFI_WRDATA_P1_slice_63;
wire   [0:0]     DFI_WRDATA_P2_slice_0;
wire   [32:32]   DFI_WRDATA_P2_slice_1;
wire   [1:1]     DFI_WRDATA_P2_slice_2;
wire   [33:33]   DFI_WRDATA_P2_slice_3;
wire   [2:2]     DFI_WRDATA_P2_slice_4;
wire   [34:34]   DFI_WRDATA_P2_slice_5;
wire   [3:3]     DFI_WRDATA_P2_slice_6;
wire   [35:35]   DFI_WRDATA_P2_slice_7;
wire   [4:4]     DFI_WRDATA_P2_slice_8;
wire   [36:36]   DFI_WRDATA_P2_slice_9;
wire   [5:5]     DFI_WRDATA_P2_slice_10;
wire   [37:37]   DFI_WRDATA_P2_slice_11;
wire   [6:6]     DFI_WRDATA_P2_slice_12;
wire   [38:38]   DFI_WRDATA_P2_slice_13;
wire   [7:7]     DFI_WRDATA_P2_slice_14;
wire   [39:39]   DFI_WRDATA_P2_slice_15;
wire   [8:8]     DFI_WRDATA_P2_slice_16;
wire   [40:40]   DFI_WRDATA_P2_slice_17;
wire   [9:9]     DFI_WRDATA_P2_slice_18;
wire   [41:41]   DFI_WRDATA_P2_slice_19;
wire   [10:10]   DFI_WRDATA_P2_slice_20;
wire   [42:42]   DFI_WRDATA_P2_slice_21;
wire   [11:11]   DFI_WRDATA_P2_slice_22;
wire   [43:43]   DFI_WRDATA_P2_slice_23;
wire   [12:12]   DFI_WRDATA_P2_slice_24;
wire   [44:44]   DFI_WRDATA_P2_slice_25;
wire   [13:13]   DFI_WRDATA_P2_slice_26;
wire   [45:45]   DFI_WRDATA_P2_slice_27;
wire   [14:14]   DFI_WRDATA_P2_slice_28;
wire   [46:46]   DFI_WRDATA_P2_slice_29;
wire   [15:15]   DFI_WRDATA_P2_slice_30;
wire   [47:47]   DFI_WRDATA_P2_slice_31;
wire   [16:16]   DFI_WRDATA_P2_slice_32;
wire   [48:48]   DFI_WRDATA_P2_slice_33;
wire   [17:17]   DFI_WRDATA_P2_slice_34;
wire   [49:49]   DFI_WRDATA_P2_slice_35;
wire   [18:18]   DFI_WRDATA_P2_slice_36;
wire   [50:50]   DFI_WRDATA_P2_slice_37;
wire   [19:19]   DFI_WRDATA_P2_slice_38;
wire   [51:51]   DFI_WRDATA_P2_slice_39;
wire   [20:20]   DFI_WRDATA_P2_slice_40;
wire   [52:52]   DFI_WRDATA_P2_slice_41;
wire   [21:21]   DFI_WRDATA_P2_slice_42;
wire   [53:53]   DFI_WRDATA_P2_slice_43;
wire   [22:22]   DFI_WRDATA_P2_slice_44;
wire   [54:54]   DFI_WRDATA_P2_slice_45;
wire   [23:23]   DFI_WRDATA_P2_slice_46;
wire   [55:55]   DFI_WRDATA_P2_slice_47;
wire   [24:24]   DFI_WRDATA_P2_slice_48;
wire   [56:56]   DFI_WRDATA_P2_slice_49;
wire   [25:25]   DFI_WRDATA_P2_slice_50;
wire   [57:57]   DFI_WRDATA_P2_slice_51;
wire   [26:26]   DFI_WRDATA_P2_slice_52;
wire   [58:58]   DFI_WRDATA_P2_slice_53;
wire   [27:27]   DFI_WRDATA_P2_slice_54;
wire   [59:59]   DFI_WRDATA_P2_slice_55;
wire   [28:28]   DFI_WRDATA_P2_slice_56;
wire   [60:60]   DFI_WRDATA_P2_slice_57;
wire   [29:29]   DFI_WRDATA_P2_slice_58;
wire   [61:61]   DFI_WRDATA_P2_slice_59;
wire   [30:30]   DFI_WRDATA_P2_slice_60;
wire   [62:62]   DFI_WRDATA_P2_slice_61;
wire   [31:31]   DFI_WRDATA_P2_slice_62;
wire   [63:63]   DFI_WRDATA_P2_slice_63;
wire   [0:0]     DFI_WRDATA_P3_slice_0;
wire   [32:32]   DFI_WRDATA_P3_slice_1;
wire   [1:1]     DFI_WRDATA_P3_slice_2;
wire   [33:33]   DFI_WRDATA_P3_slice_3;
wire   [2:2]     DFI_WRDATA_P3_slice_4;
wire   [34:34]   DFI_WRDATA_P3_slice_5;
wire   [3:3]     DFI_WRDATA_P3_slice_6;
wire   [35:35]   DFI_WRDATA_P3_slice_7;
wire   [4:4]     DFI_WRDATA_P3_slice_8;
wire   [36:36]   DFI_WRDATA_P3_slice_9;
wire   [5:5]     DFI_WRDATA_P3_slice_10;
wire   [37:37]   DFI_WRDATA_P3_slice_11;
wire   [6:6]     DFI_WRDATA_P3_slice_12;
wire   [38:38]   DFI_WRDATA_P3_slice_13;
wire   [7:7]     DFI_WRDATA_P3_slice_14;
wire   [39:39]   DFI_WRDATA_P3_slice_15;
wire   [8:8]     DFI_WRDATA_P3_slice_16;
wire   [40:40]   DFI_WRDATA_P3_slice_17;
wire   [9:9]     DFI_WRDATA_P3_slice_18;
wire   [41:41]   DFI_WRDATA_P3_slice_19;
wire   [10:10]   DFI_WRDATA_P3_slice_20;
wire   [42:42]   DFI_WRDATA_P3_slice_21;
wire   [11:11]   DFI_WRDATA_P3_slice_22;
wire   [43:43]   DFI_WRDATA_P3_slice_23;
wire   [12:12]   DFI_WRDATA_P3_slice_24;
wire   [44:44]   DFI_WRDATA_P3_slice_25;
wire   [13:13]   DFI_WRDATA_P3_slice_26;
wire   [45:45]   DFI_WRDATA_P3_slice_27;
wire   [14:14]   DFI_WRDATA_P3_slice_28;
wire   [46:46]   DFI_WRDATA_P3_slice_29;
wire   [15:15]   DFI_WRDATA_P3_slice_30;
wire   [47:47]   DFI_WRDATA_P3_slice_31;
wire   [16:16]   DFI_WRDATA_P3_slice_32;
wire   [48:48]   DFI_WRDATA_P3_slice_33;
wire   [17:17]   DFI_WRDATA_P3_slice_34;
wire   [49:49]   DFI_WRDATA_P3_slice_35;
wire   [18:18]   DFI_WRDATA_P3_slice_36;
wire   [50:50]   DFI_WRDATA_P3_slice_37;
wire   [19:19]   DFI_WRDATA_P3_slice_38;
wire   [51:51]   DFI_WRDATA_P3_slice_39;
wire   [20:20]   DFI_WRDATA_P3_slice_40;
wire   [52:52]   DFI_WRDATA_P3_slice_41;
wire   [21:21]   DFI_WRDATA_P3_slice_42;
wire   [53:53]   DFI_WRDATA_P3_slice_43;
wire   [22:22]   DFI_WRDATA_P3_slice_44;
wire   [54:54]   DFI_WRDATA_P3_slice_45;
wire   [23:23]   DFI_WRDATA_P3_slice_46;
wire   [55:55]   DFI_WRDATA_P3_slice_47;
wire   [24:24]   DFI_WRDATA_P3_slice_48;
wire   [56:56]   DFI_WRDATA_P3_slice_49;
wire   [25:25]   DFI_WRDATA_P3_slice_50;
wire   [57:57]   DFI_WRDATA_P3_slice_51;
wire   [26:26]   DFI_WRDATA_P3_slice_52;
wire   [58:58]   DFI_WRDATA_P3_slice_53;
wire   [27:27]   DFI_WRDATA_P3_slice_54;
wire   [59:59]   DFI_WRDATA_P3_slice_55;
wire   [28:28]   DFI_WRDATA_P3_slice_56;
wire   [60:60]   DFI_WRDATA_P3_slice_57;
wire   [29:29]   DFI_WRDATA_P3_slice_58;
wire   [61:61]   DFI_WRDATA_P3_slice_59;
wire   [30:30]   DFI_WRDATA_P3_slice_60;
wire   [62:62]   DFI_WRDATA_P3_slice_61;
wire   [31:31]   DFI_WRDATA_P3_slice_62;
wire   [63:63]   DFI_WRDATA_P3_slice_63;
wire   [0:0]     DFI_WRLVL_CS_N;
wire             DFI_WRLVL_EN;
wire   [3:0]     DFI_WRLVL_RESP_net_0;
wire             DFI_WRLVL_STROBE;
wire             DFN1_CMD_Q;
wire   [7:0]     DLL_CODE;
wire             DLL_DLY_DIFF;
wire   [0:0]     DM_N_net_0;
wire   [0:0]     DM_N_0;
wire   [0:0]     DM_N_1;
wire   [0:0]     DM_N_2;
wire             HS_IO_CLK;
wire             HS_IO_CLK_270;
wire             IOD_A_12_EYE_MONITOR_EARLY_0;
wire             IOD_A_12_EYE_MONITOR_LATE_0;
wire   [3:3]     IOD_A_12_RX_DATA_03to3;
wire             IOD_A_12_TX_0;
wire             IOD_BCLK_TRAINING_EYE_MONITOR_EARLY_0;
wire             IOD_BCLK_TRAINING_EYE_MONITOR_LATE_0;
wire   [0:0]     IOD_BCLK_TRAINING_RX_DATA_00to0;
wire   [2:2]     IOD_BCLK_TRAINING_RX_DATA_02to2;
wire   [4:4]     IOD_BCLK_TRAINING_RX_DATA_04to4;
wire   [6:6]     IOD_BCLK_TRAINING_RX_DATA_06to6;
wire             IOD_REF_CLK_TRAINING_EYE_MONITOR_EARLY_0;
wire             IOD_REF_CLK_TRAINING_EYE_MONITOR_LATE_0;
wire   [6:6]     IOD_REF_CLK_TRAINING_RX_DATA_06to6;
wire   [0:0]     IOD_TRAINING_0_BCLK_EYE_MONITOR_CLR_FLAGS;
wire   [0:0]     IOD_TRAINING_0_CLK_SEL0to0;
wire   [1:1]     IOD_TRAINING_0_CLK_SEL1to1;
wire   [2:2]     IOD_TRAINING_0_CLK_SEL2to2;
wire   [3:3]     IOD_TRAINING_0_CLK_SEL3to3;
wire   [4:4]     IOD_TRAINING_0_CLK_SEL4to4;
wire   [5:5]     IOD_TRAINING_0_CLK_SEL5to5;
wire   [6:6]     IOD_TRAINING_0_CLK_SEL6to6;
wire   [7:7]     IOD_TRAINING_0_CLK_SEL7to7;
wire   [8:8]     IOD_TRAINING_0_CLK_SEL8to8;
wire   [9:9]     IOD_TRAINING_0_CLK_SEL9to9;
wire   [10:10]   IOD_TRAINING_0_CLK_SEL10to10;
wire   [11:11]   IOD_TRAINING_0_CLK_SEL11to11;
wire             IOD_TRAINING_0_CMD_DELAY_LINE_DIRECTION;
wire             IOD_TRAINING_0_CMD_DELAY_LINE_LOAD;
wire             IOD_TRAINING_0_CMD_DELAY_LINE_MOVE;
wire             IOD_TRAINING_0_CMD_DELAY_LINE_MOVE_TRN;
wire             IOD_TRAINING_0_CMD_EYE_MONITOR_CLR_FLAGS;
wire             IOD_TRAINING_0_CMD_OE;
wire             IOD_TRAINING_0_CMD_RESET_LANE;
wire   [0:0]     IOD_TRAINING_0_DELAY_LINE_SEL_RD0to0;
wire   [1:1]     IOD_TRAINING_0_DELAY_LINE_SEL_RD1to1;
wire   [2:2]     IOD_TRAINING_0_DELAY_LINE_SEL_RD2to2;
wire   [3:3]     IOD_TRAINING_0_DELAY_LINE_SEL_RD3to3;
wire             IOD_TRAINING_0_DFI_ACT_N_P0_OUT;
wire             IOD_TRAINING_0_DFI_ACT_N_P1_OUT;
wire             IOD_TRAINING_0_DFI_ACT_N_P2_OUT;
wire             IOD_TRAINING_0_DFI_ACT_N_P3_OUT;
wire   [0:0]     IOD_TRAINING_0_DFI_BANK_P0_OUT0to0;
wire   [1:1]     IOD_TRAINING_0_DFI_BANK_P0_OUT1to1;
wire   [0:0]     IOD_TRAINING_0_DFI_BANK_P1_OUT0to0;
wire   [1:1]     IOD_TRAINING_0_DFI_BANK_P1_OUT1to1;
wire   [0:0]     IOD_TRAINING_0_DFI_BANK_P2_OUT0to0;
wire   [1:1]     IOD_TRAINING_0_DFI_BANK_P2_OUT1to1;
wire   [0:0]     IOD_TRAINING_0_DFI_BANK_P3_OUT0to0;
wire   [1:1]     IOD_TRAINING_0_DFI_BANK_P3_OUT1to1;
wire   [0:0]     IOD_TRAINING_0_DFI_BG_P0_OUT0to0;
wire   [1:1]     IOD_TRAINING_0_DFI_BG_P0_OUT1to1;
wire   [0:0]     IOD_TRAINING_0_DFI_BG_P1_OUT0to0;
wire   [1:1]     IOD_TRAINING_0_DFI_BG_P1_OUT1to1;
wire   [0:0]     IOD_TRAINING_0_DFI_BG_P2_OUT0to0;
wire   [1:1]     IOD_TRAINING_0_DFI_BG_P2_OUT1to1;
wire   [0:0]     IOD_TRAINING_0_DFI_BG_P3_OUT0to0;
wire   [1:1]     IOD_TRAINING_0_DFI_BG_P3_OUT1to1;
wire             IOD_TRAINING_0_DFI_CAS_N_P0_OUT;
wire             IOD_TRAINING_0_DFI_CAS_N_P1_OUT;
wire             IOD_TRAINING_0_DFI_CAS_N_P2_OUT;
wire             IOD_TRAINING_0_DFI_CAS_N_P3_OUT;
wire             IOD_TRAINING_0_DFI_CKE_P0_OUT;
wire             IOD_TRAINING_0_DFI_CKE_P1_OUT;
wire             IOD_TRAINING_0_DFI_CKE_P2_OUT;
wire             IOD_TRAINING_0_DFI_CKE_P3_OUT;
wire             IOD_TRAINING_0_DFI_CS_N_P0_OUT;
wire             IOD_TRAINING_0_DFI_CS_N_P1_OUT;
wire             IOD_TRAINING_0_DFI_CS_N_P2_OUT;
wire             IOD_TRAINING_0_DFI_CS_N_P3_OUT;
wire             IOD_TRAINING_0_DFI_ODT_P0_OUT;
wire             IOD_TRAINING_0_DFI_ODT_P1_OUT;
wire             IOD_TRAINING_0_DFI_ODT_P2_OUT;
wire             IOD_TRAINING_0_DFI_ODT_P3_OUT;
wire             IOD_TRAINING_0_DFI_RAS_N_P0_OUT;
wire             IOD_TRAINING_0_DFI_RAS_N_P1_OUT;
wire             IOD_TRAINING_0_DFI_RAS_N_P2_OUT;
wire             IOD_TRAINING_0_DFI_RAS_N_P3_OUT;
wire             IOD_TRAINING_0_DFI_RESET_N_P0_OUT;
wire             IOD_TRAINING_0_DFI_RESET_N_P1_OUT;
wire             IOD_TRAINING_0_DFI_RESET_N_P2_OUT;
wire             IOD_TRAINING_0_DFI_RESET_N_P3_OUT;
wire             IOD_TRAINING_0_DFI_WE_N_P0_OUT;
wire             IOD_TRAINING_0_DFI_WE_N_P1_OUT;
wire             IOD_TRAINING_0_DFI_WE_N_P2_OUT;
wire             IOD_TRAINING_0_DFI_WE_N_P3_OUT;
wire   [0:0]     IOD_TRAINING_0_DIRECTION0to0;
wire   [1:1]     IOD_TRAINING_0_DIRECTION1to1;
wire   [2:2]     IOD_TRAINING_0_DIRECTION2to2;
wire   [3:3]     IOD_TRAINING_0_DIRECTION3to3;
wire   [4:4]     IOD_TRAINING_0_DIRECTION4to4;
wire   [5:5]     IOD_TRAINING_0_DIRECTION5to5;
wire   [6:6]     IOD_TRAINING_0_DIRECTION6to6;
wire   [7:7]     IOD_TRAINING_0_DIRECTION7to7;
wire   [8:8]     IOD_TRAINING_0_DIRECTION8to8;
wire   [9:9]     IOD_TRAINING_0_DIRECTION9to9;
wire   [10:10]   IOD_TRAINING_0_DIRECTION10to10;
wire   [11:11]   IOD_TRAINING_0_DIRECTION11to11;
wire   [12:12]   IOD_TRAINING_0_DIRECTION12to12;
wire   [13:13]   IOD_TRAINING_0_DIRECTION13to13;
wire   [14:14]   IOD_TRAINING_0_DIRECTION14to14;
wire   [15:15]   IOD_TRAINING_0_DIRECTION15to15;
wire   [16:16]   IOD_TRAINING_0_DIRECTION16to16;
wire   [17:17]   IOD_TRAINING_0_DIRECTION17to17;
wire   [18:18]   IOD_TRAINING_0_DIRECTION18to18;
wire   [19:19]   IOD_TRAINING_0_DIRECTION19to19;
wire   [20:20]   IOD_TRAINING_0_DIRECTION20to20;
wire   [21:21]   IOD_TRAINING_0_DIRECTION21to21;
wire   [22:22]   IOD_TRAINING_0_DIRECTION22to22;
wire   [23:23]   IOD_TRAINING_0_DIRECTION23to23;
wire   [24:24]   IOD_TRAINING_0_DIRECTION24to24;
wire   [25:25]   IOD_TRAINING_0_DIRECTION25to25;
wire   [26:26]   IOD_TRAINING_0_DIRECTION26to26;
wire   [27:27]   IOD_TRAINING_0_DIRECTION27to27;
wire   [28:28]   IOD_TRAINING_0_DIRECTION28to28;
wire   [29:29]   IOD_TRAINING_0_DIRECTION29to29;
wire   [30:30]   IOD_TRAINING_0_DIRECTION30to30;
wire   [31:31]   IOD_TRAINING_0_DIRECTION31to31;
wire   [32:32]   IOD_TRAINING_0_DIRECTION32to32;
wire   [33:33]   IOD_TRAINING_0_DIRECTION33to33;
wire   [34:34]   IOD_TRAINING_0_DIRECTION34to34;
wire   [35:35]   IOD_TRAINING_0_DIRECTION35to35;
wire   [0:0]     IOD_TRAINING_0_DM_OE_P00to0;
wire   [1:1]     IOD_TRAINING_0_DM_OE_P01to1;
wire   [2:2]     IOD_TRAINING_0_DM_OE_P02to2;
wire   [3:3]     IOD_TRAINING_0_DM_OE_P03to3;
wire   [0:0]     IOD_TRAINING_0_DM_OE_P10to0;
wire   [1:1]     IOD_TRAINING_0_DM_OE_P11to1;
wire   [2:2]     IOD_TRAINING_0_DM_OE_P12to2;
wire   [3:3]     IOD_TRAINING_0_DM_OE_P13to3;
wire   [0:0]     IOD_TRAINING_0_DM_OE_P20to0;
wire   [1:1]     IOD_TRAINING_0_DM_OE_P21to1;
wire   [2:2]     IOD_TRAINING_0_DM_OE_P22to2;
wire   [3:3]     IOD_TRAINING_0_DM_OE_P23to3;
wire   [0:0]     IOD_TRAINING_0_DM_OE_P30to0;
wire   [1:1]     IOD_TRAINING_0_DM_OE_P31to1;
wire   [2:2]     IOD_TRAINING_0_DM_OE_P32to2;
wire   [3:3]     IOD_TRAINING_0_DM_OE_P33to3;
wire   [0:0]     IOD_TRAINING_0_DQS_OE_P00to0;
wire   [1:1]     IOD_TRAINING_0_DQS_OE_P01to1;
wire   [2:2]     IOD_TRAINING_0_DQS_OE_P02to2;
wire   [3:3]     IOD_TRAINING_0_DQS_OE_P03to3;
wire   [0:0]     IOD_TRAINING_0_DQS_OE_P10to0;
wire   [1:1]     IOD_TRAINING_0_DQS_OE_P11to1;
wire   [2:2]     IOD_TRAINING_0_DQS_OE_P12to2;
wire   [3:3]     IOD_TRAINING_0_DQS_OE_P13to3;
wire   [0:0]     IOD_TRAINING_0_DQS_OE_P20to0;
wire   [1:1]     IOD_TRAINING_0_DQS_OE_P21to1;
wire   [2:2]     IOD_TRAINING_0_DQS_OE_P22to2;
wire   [3:3]     IOD_TRAINING_0_DQS_OE_P23to3;
wire   [0:0]     IOD_TRAINING_0_DQS_OE_P30to0;
wire   [1:1]     IOD_TRAINING_0_DQS_OE_P31to1;
wire   [2:2]     IOD_TRAINING_0_DQS_OE_P32to2;
wire   [3:3]     IOD_TRAINING_0_DQS_OE_P33to3;
wire   [0:0]     IOD_TRAINING_0_DQSW270_DELAY_LINE_DIRECTION0to0;
wire   [1:1]     IOD_TRAINING_0_DQSW270_DELAY_LINE_DIRECTION1to1;
wire   [2:2]     IOD_TRAINING_0_DQSW270_DELAY_LINE_DIRECTION2to2;
wire   [3:3]     IOD_TRAINING_0_DQSW270_DELAY_LINE_DIRECTION3to3;
wire   [0:0]     IOD_TRAINING_0_DQSW270_DELAY_LINE_LOAD0to0;
wire   [1:1]     IOD_TRAINING_0_DQSW270_DELAY_LINE_LOAD1to1;
wire   [2:2]     IOD_TRAINING_0_DQSW270_DELAY_LINE_LOAD2to2;
wire   [3:3]     IOD_TRAINING_0_DQSW270_DELAY_LINE_LOAD3to3;
wire   [0:0]     IOD_TRAINING_0_DQSW270_DELAY_LINE_MOVE0to0;
wire   [1:1]     IOD_TRAINING_0_DQSW270_DELAY_LINE_MOVE1to1;
wire   [2:2]     IOD_TRAINING_0_DQSW270_DELAY_LINE_MOVE2to2;
wire   [3:3]     IOD_TRAINING_0_DQSW270_DELAY_LINE_MOVE3to3;
wire   [0:0]     IOD_TRAINING_0_DQSW270_EYE_MONITOR_CLR_FLAGS0to0;
wire   [1:1]     IOD_TRAINING_0_DQSW270_EYE_MONITOR_CLR_FLAGS1to1;
wire   [2:2]     IOD_TRAINING_0_DQSW270_EYE_MONITOR_CLR_FLAGS2to2;
wire   [3:3]     IOD_TRAINING_0_DQSW270_EYE_MONITOR_CLR_FLAGS3to3;
wire   [0:0]     IOD_TRAINING_0_DQSW_DELAY_LINE_DIRECTION0to0;
wire   [1:1]     IOD_TRAINING_0_DQSW_DELAY_LINE_DIRECTION1to1;
wire   [2:2]     IOD_TRAINING_0_DQSW_DELAY_LINE_DIRECTION2to2;
wire   [3:3]     IOD_TRAINING_0_DQSW_DELAY_LINE_DIRECTION3to3;
wire   [0:0]     IOD_TRAINING_0_DQSW_DELAY_LINE_LOAD0to0;
wire   [1:1]     IOD_TRAINING_0_DQSW_DELAY_LINE_LOAD1to1;
wire   [2:2]     IOD_TRAINING_0_DQSW_DELAY_LINE_LOAD2to2;
wire   [3:3]     IOD_TRAINING_0_DQSW_DELAY_LINE_LOAD3to3;
wire   [0:0]     IOD_TRAINING_0_DQSW_DELAY_LINE_MOVE0to0;
wire   [1:1]     IOD_TRAINING_0_DQSW_DELAY_LINE_MOVE1to1;
wire   [2:2]     IOD_TRAINING_0_DQSW_DELAY_LINE_MOVE2to2;
wire   [3:3]     IOD_TRAINING_0_DQSW_DELAY_LINE_MOVE3to3;
wire   [0:0]     IOD_TRAINING_0_DQSW_EYE_MONITOR_CLR_FLAGS0to0;
wire   [1:1]     IOD_TRAINING_0_DQSW_EYE_MONITOR_CLR_FLAGS1to1;
wire   [2:2]     IOD_TRAINING_0_DQSW_EYE_MONITOR_CLR_FLAGS2to2;
wire   [3:3]     IOD_TRAINING_0_DQSW_EYE_MONITOR_CLR_FLAGS3to3;
wire   [7:0]     IOD_TRAINING_0_DQSW_SELA7to0;
wire   [15:8]    IOD_TRAINING_0_DQSW_SELA15to8;
wire   [23:16]   IOD_TRAINING_0_DQSW_SELA23to16;
wire   [31:24]   IOD_TRAINING_0_DQSW_SELA31to24;
wire   [0:0]     IOD_TRAINING_0_INIT_PAUSE0to0;
wire   [1:1]     IOD_TRAINING_0_INIT_PAUSE1to1;
wire   [2:2]     IOD_TRAINING_0_INIT_PAUSE2to2;
wire   [3:3]     IOD_TRAINING_0_INIT_PAUSE3to3;
wire   [0:0]     IOD_TRAINING_0_IOG_ADDRESS_P00to0;
wire   [1:1]     IOD_TRAINING_0_IOG_ADDRESS_P01to1;
wire   [2:2]     IOD_TRAINING_0_IOG_ADDRESS_P02to2;
wire   [3:3]     IOD_TRAINING_0_IOG_ADDRESS_P03to3;
wire   [4:4]     IOD_TRAINING_0_IOG_ADDRESS_P04to4;
wire   [5:5]     IOD_TRAINING_0_IOG_ADDRESS_P05to5;
wire   [6:6]     IOD_TRAINING_0_IOG_ADDRESS_P06to6;
wire   [7:7]     IOD_TRAINING_0_IOG_ADDRESS_P07to7;
wire   [8:8]     IOD_TRAINING_0_IOG_ADDRESS_P08to8;
wire   [9:9]     IOD_TRAINING_0_IOG_ADDRESS_P09to9;
wire   [0:0]     IOD_TRAINING_0_IOG_ADDRESS_P10to0;
wire   [10:10]   IOD_TRAINING_0_IOG_ADDRESS_P010to10;
wire   [1:1]     IOD_TRAINING_0_IOG_ADDRESS_P11to1;
wire   [11:11]   IOD_TRAINING_0_IOG_ADDRESS_P011to11;
wire   [2:2]     IOD_TRAINING_0_IOG_ADDRESS_P12to2;
wire   [12:12]   IOD_TRAINING_0_IOG_ADDRESS_P012to12;
wire   [3:3]     IOD_TRAINING_0_IOG_ADDRESS_P13to3;
wire   [13:13]   IOD_TRAINING_0_IOG_ADDRESS_P013to13;
wire   [4:4]     IOD_TRAINING_0_IOG_ADDRESS_P14to4;
wire   [5:5]     IOD_TRAINING_0_IOG_ADDRESS_P15to5;
wire   [6:6]     IOD_TRAINING_0_IOG_ADDRESS_P16to6;
wire   [7:7]     IOD_TRAINING_0_IOG_ADDRESS_P17to7;
wire   [8:8]     IOD_TRAINING_0_IOG_ADDRESS_P18to8;
wire   [9:9]     IOD_TRAINING_0_IOG_ADDRESS_P19to9;
wire   [0:0]     IOD_TRAINING_0_IOG_ADDRESS_P20to0;
wire   [1:1]     IOD_TRAINING_0_IOG_ADDRESS_P21to1;
wire   [2:2]     IOD_TRAINING_0_IOG_ADDRESS_P22to2;
wire   [3:3]     IOD_TRAINING_0_IOG_ADDRESS_P23to3;
wire   [4:4]     IOD_TRAINING_0_IOG_ADDRESS_P24to4;
wire   [5:5]     IOD_TRAINING_0_IOG_ADDRESS_P25to5;
wire   [6:6]     IOD_TRAINING_0_IOG_ADDRESS_P26to6;
wire   [7:7]     IOD_TRAINING_0_IOG_ADDRESS_P27to7;
wire   [8:8]     IOD_TRAINING_0_IOG_ADDRESS_P28to8;
wire   [9:9]     IOD_TRAINING_0_IOG_ADDRESS_P29to9;
wire   [0:0]     IOD_TRAINING_0_IOG_ADDRESS_P30to0;
wire   [1:1]     IOD_TRAINING_0_IOG_ADDRESS_P31to1;
wire   [2:2]     IOD_TRAINING_0_IOG_ADDRESS_P32to2;
wire   [3:3]     IOD_TRAINING_0_IOG_ADDRESS_P33to3;
wire   [4:4]     IOD_TRAINING_0_IOG_ADDRESS_P34to4;
wire   [5:5]     IOD_TRAINING_0_IOG_ADDRESS_P35to5;
wire   [6:6]     IOD_TRAINING_0_IOG_ADDRESS_P36to6;
wire   [7:7]     IOD_TRAINING_0_IOG_ADDRESS_P37to7;
wire   [8:8]     IOD_TRAINING_0_IOG_ADDRESS_P38to8;
wire   [9:9]     IOD_TRAINING_0_IOG_ADDRESS_P39to9;
wire   [10:10]   IOD_TRAINING_0_IOG_ADDRESS_P110to10;
wire   [11:11]   IOD_TRAINING_0_IOG_ADDRESS_P111to11;
wire   [12:12]   IOD_TRAINING_0_IOG_ADDRESS_P112to12;
wire   [13:13]   IOD_TRAINING_0_IOG_ADDRESS_P113to13;
wire   [10:10]   IOD_TRAINING_0_IOG_ADDRESS_P210to10;
wire   [11:11]   IOD_TRAINING_0_IOG_ADDRESS_P211to11;
wire   [12:12]   IOD_TRAINING_0_IOG_ADDRESS_P212to12;
wire   [13:13]   IOD_TRAINING_0_IOG_ADDRESS_P213to13;
wire   [10:10]   IOD_TRAINING_0_IOG_ADDRESS_P310to10;
wire   [11:11]   IOD_TRAINING_0_IOG_ADDRESS_P311to11;
wire   [12:12]   IOD_TRAINING_0_IOG_ADDRESS_P312to12;
wire   [13:13]   IOD_TRAINING_0_IOG_ADDRESS_P313to13;
wire   [0:0]     IOD_TRAINING_0_IOG_DM_TXDATA_OUT0to0;
wire   [1:1]     IOD_TRAINING_0_IOG_DM_TXDATA_OUT1to1;
wire   [2:2]     IOD_TRAINING_0_IOG_DM_TXDATA_OUT2to2;
wire   [3:3]     IOD_TRAINING_0_IOG_DM_TXDATA_OUT3to3;
wire   [4:4]     IOD_TRAINING_0_IOG_DM_TXDATA_OUT4to4;
wire   [5:5]     IOD_TRAINING_0_IOG_DM_TXDATA_OUT5to5;
wire   [6:6]     IOD_TRAINING_0_IOG_DM_TXDATA_OUT6to6;
wire   [7:7]     IOD_TRAINING_0_IOG_DM_TXDATA_OUT7to7;
wire   [8:8]     IOD_TRAINING_0_IOG_DM_TXDATA_OUT8to8;
wire   [9:9]     IOD_TRAINING_0_IOG_DM_TXDATA_OUT9to9;
wire   [10:10]   IOD_TRAINING_0_IOG_DM_TXDATA_OUT10to10;
wire   [11:11]   IOD_TRAINING_0_IOG_DM_TXDATA_OUT11to11;
wire   [12:12]   IOD_TRAINING_0_IOG_DM_TXDATA_OUT12to12;
wire   [13:13]   IOD_TRAINING_0_IOG_DM_TXDATA_OUT13to13;
wire   [14:14]   IOD_TRAINING_0_IOG_DM_TXDATA_OUT14to14;
wire   [15:15]   IOD_TRAINING_0_IOG_DM_TXDATA_OUT15to15;
wire   [16:16]   IOD_TRAINING_0_IOG_DM_TXDATA_OUT16to16;
wire   [17:17]   IOD_TRAINING_0_IOG_DM_TXDATA_OUT17to17;
wire   [18:18]   IOD_TRAINING_0_IOG_DM_TXDATA_OUT18to18;
wire   [19:19]   IOD_TRAINING_0_IOG_DM_TXDATA_OUT19to19;
wire   [20:20]   IOD_TRAINING_0_IOG_DM_TXDATA_OUT20to20;
wire   [21:21]   IOD_TRAINING_0_IOG_DM_TXDATA_OUT21to21;
wire   [22:22]   IOD_TRAINING_0_IOG_DM_TXDATA_OUT22to22;
wire   [23:23]   IOD_TRAINING_0_IOG_DM_TXDATA_OUT23to23;
wire   [24:24]   IOD_TRAINING_0_IOG_DM_TXDATA_OUT24to24;
wire   [25:25]   IOD_TRAINING_0_IOG_DM_TXDATA_OUT25to25;
wire   [26:26]   IOD_TRAINING_0_IOG_DM_TXDATA_OUT26to26;
wire   [27:27]   IOD_TRAINING_0_IOG_DM_TXDATA_OUT27to27;
wire   [28:28]   IOD_TRAINING_0_IOG_DM_TXDATA_OUT28to28;
wire   [29:29]   IOD_TRAINING_0_IOG_DM_TXDATA_OUT29to29;
wire   [30:30]   IOD_TRAINING_0_IOG_DM_TXDATA_OUT30to30;
wire   [31:31]   IOD_TRAINING_0_IOG_DM_TXDATA_OUT31to31;
wire   [0:0]     IOD_TRAINING_0_IOG_DQ_TXDATA_OUT0to0;
wire   [1:1]     IOD_TRAINING_0_IOG_DQ_TXDATA_OUT1to1;
wire   [2:2]     IOD_TRAINING_0_IOG_DQ_TXDATA_OUT2to2;
wire   [3:3]     IOD_TRAINING_0_IOG_DQ_TXDATA_OUT3to3;
wire   [4:4]     IOD_TRAINING_0_IOG_DQ_TXDATA_OUT4to4;
wire   [5:5]     IOD_TRAINING_0_IOG_DQ_TXDATA_OUT5to5;
wire   [6:6]     IOD_TRAINING_0_IOG_DQ_TXDATA_OUT6to6;
wire   [7:7]     IOD_TRAINING_0_IOG_DQ_TXDATA_OUT7to7;
wire   [8:8]     IOD_TRAINING_0_IOG_DQ_TXDATA_OUT8to8;
wire   [9:9]     IOD_TRAINING_0_IOG_DQ_TXDATA_OUT9to9;
wire   [10:10]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT10to10;
wire   [11:11]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT11to11;
wire   [12:12]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT12to12;
wire   [13:13]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT13to13;
wire   [14:14]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT14to14;
wire   [15:15]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT15to15;
wire   [16:16]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT16to16;
wire   [17:17]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT17to17;
wire   [18:18]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT18to18;
wire   [19:19]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT19to19;
wire   [20:20]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT20to20;
wire   [21:21]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT21to21;
wire   [22:22]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT22to22;
wire   [23:23]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT23to23;
wire   [24:24]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT24to24;
wire   [25:25]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT25to25;
wire   [26:26]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT26to26;
wire   [27:27]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT27to27;
wire   [28:28]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT28to28;
wire   [29:29]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT29to29;
wire   [30:30]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT30to30;
wire   [31:31]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT31to31;
wire   [32:32]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT32to32;
wire   [33:33]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT33to33;
wire   [34:34]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT34to34;
wire   [35:35]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT35to35;
wire   [36:36]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT36to36;
wire   [37:37]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT37to37;
wire   [38:38]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT38to38;
wire   [39:39]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT39to39;
wire   [40:40]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT40to40;
wire   [41:41]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT41to41;
wire   [42:42]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT42to42;
wire   [43:43]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT43to43;
wire   [44:44]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT44to44;
wire   [45:45]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT45to45;
wire   [46:46]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT46to46;
wire   [47:47]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT47to47;
wire   [48:48]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT48to48;
wire   [49:49]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT49to49;
wire   [50:50]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT50to50;
wire   [51:51]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT51to51;
wire   [52:52]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT52to52;
wire   [53:53]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT53to53;
wire   [54:54]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT54to54;
wire   [55:55]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT55to55;
wire   [56:56]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT56to56;
wire   [57:57]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT57to57;
wire   [58:58]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT58to58;
wire   [59:59]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT59to59;
wire   [60:60]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT60to60;
wire   [61:61]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT61to61;
wire   [62:62]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT62to62;
wire   [63:63]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT63to63;
wire   [64:64]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT64to64;
wire   [65:65]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT65to65;
wire   [66:66]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT66to66;
wire   [67:67]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT67to67;
wire   [68:68]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT68to68;
wire   [69:69]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT69to69;
wire   [70:70]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT70to70;
wire   [71:71]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT71to71;
wire   [72:72]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT72to72;
wire   [73:73]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT73to73;
wire   [74:74]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT74to74;
wire   [75:75]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT75to75;
wire   [76:76]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT76to76;
wire   [77:77]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT77to77;
wire   [78:78]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT78to78;
wire   [79:79]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT79to79;
wire   [80:80]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT80to80;
wire   [81:81]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT81to81;
wire   [82:82]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT82to82;
wire   [83:83]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT83to83;
wire   [84:84]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT84to84;
wire   [85:85]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT85to85;
wire   [86:86]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT86to86;
wire   [87:87]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT87to87;
wire   [88:88]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT88to88;
wire   [89:89]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT89to89;
wire   [90:90]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT90to90;
wire   [91:91]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT91to91;
wire   [92:92]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT92to92;
wire   [93:93]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT93to93;
wire   [94:94]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT94to94;
wire   [95:95]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT95to95;
wire   [96:96]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT96to96;
wire   [97:97]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT97to97;
wire   [98:98]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT98to98;
wire   [99:99]   IOD_TRAINING_0_IOG_DQ_TXDATA_OUT99to99;
wire   [100:100] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT100to100;
wire   [101:101] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT101to101;
wire   [102:102] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT102to102;
wire   [103:103] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT103to103;
wire   [104:104] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT104to104;
wire   [105:105] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT105to105;
wire   [106:106] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT106to106;
wire   [107:107] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT107to107;
wire   [108:108] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT108to108;
wire   [109:109] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT109to109;
wire   [110:110] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT110to110;
wire   [111:111] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT111to111;
wire   [112:112] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT112to112;
wire   [113:113] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT113to113;
wire   [114:114] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT114to114;
wire   [115:115] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT115to115;
wire   [116:116] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT116to116;
wire   [117:117] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT117to117;
wire   [118:118] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT118to118;
wire   [119:119] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT119to119;
wire   [120:120] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT120to120;
wire   [121:121] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT121to121;
wire   [122:122] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT122to122;
wire   [123:123] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT123to123;
wire   [124:124] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT124to124;
wire   [125:125] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT125to125;
wire   [126:126] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT126to126;
wire   [127:127] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT127to127;
wire   [128:128] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT128to128;
wire   [129:129] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT129to129;
wire   [130:130] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT130to130;
wire   [131:131] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT131to131;
wire   [132:132] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT132to132;
wire   [133:133] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT133to133;
wire   [134:134] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT134to134;
wire   [135:135] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT135to135;
wire   [136:136] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT136to136;
wire   [137:137] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT137to137;
wire   [138:138] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT138to138;
wire   [139:139] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT139to139;
wire   [140:140] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT140to140;
wire   [141:141] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT141to141;
wire   [142:142] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT142to142;
wire   [143:143] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT143to143;
wire   [144:144] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT144to144;
wire   [145:145] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT145to145;
wire   [146:146] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT146to146;
wire   [147:147] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT147to147;
wire   [148:148] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT148to148;
wire   [149:149] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT149to149;
wire   [150:150] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT150to150;
wire   [151:151] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT151to151;
wire   [152:152] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT152to152;
wire   [153:153] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT153to153;
wire   [154:154] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT154to154;
wire   [155:155] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT155to155;
wire   [156:156] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT156to156;
wire   [157:157] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT157to157;
wire   [158:158] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT158to158;
wire   [159:159] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT159to159;
wire   [160:160] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT160to160;
wire   [161:161] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT161to161;
wire   [162:162] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT162to162;
wire   [163:163] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT163to163;
wire   [164:164] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT164to164;
wire   [165:165] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT165to165;
wire   [166:166] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT166to166;
wire   [167:167] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT167to167;
wire   [168:168] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT168to168;
wire   [169:169] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT169to169;
wire   [170:170] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT170to170;
wire   [171:171] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT171to171;
wire   [172:172] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT172to172;
wire   [173:173] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT173to173;
wire   [174:174] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT174to174;
wire   [175:175] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT175to175;
wire   [176:176] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT176to176;
wire   [177:177] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT177to177;
wire   [178:178] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT178to178;
wire   [179:179] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT179to179;
wire   [180:180] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT180to180;
wire   [181:181] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT181to181;
wire   [182:182] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT182to182;
wire   [183:183] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT183to183;
wire   [184:184] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT184to184;
wire   [185:185] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT185to185;
wire   [186:186] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT186to186;
wire   [187:187] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT187to187;
wire   [188:188] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT188to188;
wire   [189:189] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT189to189;
wire   [190:190] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT190to190;
wire   [191:191] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT191to191;
wire   [192:192] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT192to192;
wire   [193:193] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT193to193;
wire   [194:194] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT194to194;
wire   [195:195] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT195to195;
wire   [196:196] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT196to196;
wire   [197:197] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT197to197;
wire   [198:198] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT198to198;
wire   [199:199] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT199to199;
wire   [200:200] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT200to200;
wire   [201:201] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT201to201;
wire   [202:202] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT202to202;
wire   [203:203] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT203to203;
wire   [204:204] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT204to204;
wire   [205:205] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT205to205;
wire   [206:206] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT206to206;
wire   [207:207] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT207to207;
wire   [208:208] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT208to208;
wire   [209:209] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT209to209;
wire   [210:210] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT210to210;
wire   [211:211] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT211to211;
wire   [212:212] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT212to212;
wire   [213:213] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT213to213;
wire   [214:214] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT214to214;
wire   [215:215] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT215to215;
wire   [216:216] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT216to216;
wire   [217:217] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT217to217;
wire   [218:218] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT218to218;
wire   [219:219] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT219to219;
wire   [220:220] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT220to220;
wire   [221:221] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT221to221;
wire   [222:222] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT222to222;
wire   [223:223] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT223to223;
wire   [224:224] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT224to224;
wire   [225:225] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT225to225;
wire   [226:226] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT226to226;
wire   [227:227] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT227to227;
wire   [228:228] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT228to228;
wire   [229:229] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT229to229;
wire   [230:230] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT230to230;
wire   [231:231] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT231to231;
wire   [232:232] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT232to232;
wire   [233:233] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT233to233;
wire   [234:234] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT234to234;
wire   [235:235] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT235to235;
wire   [236:236] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT236to236;
wire   [237:237] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT237to237;
wire   [238:238] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT238to238;
wire   [239:239] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT239to239;
wire   [240:240] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT240to240;
wire   [241:241] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT241to241;
wire   [242:242] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT242to242;
wire   [243:243] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT243to243;
wire   [244:244] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT244to244;
wire   [245:245] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT245to245;
wire   [246:246] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT246to246;
wire   [247:247] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT247to247;
wire   [248:248] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT248to248;
wire   [249:249] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT249to249;
wire   [250:250] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT250to250;
wire   [251:251] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT251to251;
wire   [252:252] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT252to252;
wire   [253:253] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT253to253;
wire   [254:254] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT254to254;
wire   [255:255] IOD_TRAINING_0_IOG_DQ_TXDATA_OUT255to255;
wire   [0:0]     IOD_TRAINING_0_IOG_OE_P00to0;
wire   [1:1]     IOD_TRAINING_0_IOG_OE_P01to1;
wire   [2:2]     IOD_TRAINING_0_IOG_OE_P02to2;
wire   [3:3]     IOD_TRAINING_0_IOG_OE_P03to3;
wire   [0:0]     IOD_TRAINING_0_IOG_OE_P10to0;
wire   [1:1]     IOD_TRAINING_0_IOG_OE_P11to1;
wire   [2:2]     IOD_TRAINING_0_IOG_OE_P12to2;
wire   [3:3]     IOD_TRAINING_0_IOG_OE_P13to3;
wire   [0:0]     IOD_TRAINING_0_IOG_OE_P20to0;
wire   [1:1]     IOD_TRAINING_0_IOG_OE_P21to1;
wire   [2:2]     IOD_TRAINING_0_IOG_OE_P22to2;
wire   [3:3]     IOD_TRAINING_0_IOG_OE_P23to3;
wire   [0:0]     IOD_TRAINING_0_IOG_OE_P30to0;
wire   [1:1]     IOD_TRAINING_0_IOG_OE_P31to1;
wire   [2:2]     IOD_TRAINING_0_IOG_OE_P32to2;
wire   [3:3]     IOD_TRAINING_0_IOG_OE_P33to3;
wire   [0:0]     IOD_TRAINING_0_IOG_RDDATA_EN_P0_N0to0;
wire   [1:1]     IOD_TRAINING_0_IOG_RDDATA_EN_P0_N1to1;
wire   [2:2]     IOD_TRAINING_0_IOG_RDDATA_EN_P0_N2to2;
wire   [3:3]     IOD_TRAINING_0_IOG_RDDATA_EN_P0_N3to3;
wire   [0:0]     IOD_TRAINING_0_IOG_RDDATA_EN_P0_P0to0;
wire   [1:1]     IOD_TRAINING_0_IOG_RDDATA_EN_P0_P1to1;
wire   [2:2]     IOD_TRAINING_0_IOG_RDDATA_EN_P0_P2to2;
wire   [3:3]     IOD_TRAINING_0_IOG_RDDATA_EN_P0_P3to3;
wire   [0:0]     IOD_TRAINING_0_IOG_RDDATA_EN_P1_N0to0;
wire   [1:1]     IOD_TRAINING_0_IOG_RDDATA_EN_P1_N1to1;
wire   [2:2]     IOD_TRAINING_0_IOG_RDDATA_EN_P1_N2to2;
wire   [3:3]     IOD_TRAINING_0_IOG_RDDATA_EN_P1_N3to3;
wire   [0:0]     IOD_TRAINING_0_IOG_RDDATA_EN_P1_P0to0;
wire   [1:1]     IOD_TRAINING_0_IOG_RDDATA_EN_P1_P1to1;
wire   [2:2]     IOD_TRAINING_0_IOG_RDDATA_EN_P1_P2to2;
wire   [3:3]     IOD_TRAINING_0_IOG_RDDATA_EN_P1_P3to3;
wire   [0:0]     IOD_TRAINING_0_IOG_RDDATA_EN_P2_N0to0;
wire   [1:1]     IOD_TRAINING_0_IOG_RDDATA_EN_P2_N1to1;
wire   [2:2]     IOD_TRAINING_0_IOG_RDDATA_EN_P2_N2to2;
wire   [3:3]     IOD_TRAINING_0_IOG_RDDATA_EN_P2_N3to3;
wire   [0:0]     IOD_TRAINING_0_IOG_RDDATA_EN_P2_P0to0;
wire   [1:1]     IOD_TRAINING_0_IOG_RDDATA_EN_P2_P1to1;
wire   [2:2]     IOD_TRAINING_0_IOG_RDDATA_EN_P2_P2to2;
wire   [3:3]     IOD_TRAINING_0_IOG_RDDATA_EN_P2_P3to3;
wire   [0:0]     IOD_TRAINING_0_IOG_RDDATA_EN_P3_N0to0;
wire   [1:1]     IOD_TRAINING_0_IOG_RDDATA_EN_P3_N1to1;
wire   [2:2]     IOD_TRAINING_0_IOG_RDDATA_EN_P3_N2to2;
wire   [3:3]     IOD_TRAINING_0_IOG_RDDATA_EN_P3_N3to3;
wire   [0:0]     IOD_TRAINING_0_IOG_RDDATA_EN_P3_P0to0;
wire   [1:1]     IOD_TRAINING_0_IOG_RDDATA_EN_P3_P1to1;
wire   [2:2]     IOD_TRAINING_0_IOG_RDDATA_EN_P3_P2to2;
wire   [3:3]     IOD_TRAINING_0_IOG_RDDATA_EN_P3_P3to3;
wire   [0:0]     IOD_TRAINING_0_LOAD0to0;
wire   [1:1]     IOD_TRAINING_0_LOAD1to1;
wire   [2:2]     IOD_TRAINING_0_LOAD2to2;
wire   [3:3]     IOD_TRAINING_0_LOAD3to3;
wire   [4:4]     IOD_TRAINING_0_LOAD4to4;
wire   [5:5]     IOD_TRAINING_0_LOAD5to5;
wire   [6:6]     IOD_TRAINING_0_LOAD6to6;
wire   [7:7]     IOD_TRAINING_0_LOAD7to7;
wire   [8:8]     IOD_TRAINING_0_LOAD8to8;
wire   [9:9]     IOD_TRAINING_0_LOAD9to9;
wire   [10:10]   IOD_TRAINING_0_LOAD10to10;
wire   [11:11]   IOD_TRAINING_0_LOAD11to11;
wire   [12:12]   IOD_TRAINING_0_LOAD12to12;
wire   [13:13]   IOD_TRAINING_0_LOAD13to13;
wire   [14:14]   IOD_TRAINING_0_LOAD14to14;
wire   [15:15]   IOD_TRAINING_0_LOAD15to15;
wire   [16:16]   IOD_TRAINING_0_LOAD16to16;
wire   [17:17]   IOD_TRAINING_0_LOAD17to17;
wire   [18:18]   IOD_TRAINING_0_LOAD18to18;
wire   [19:19]   IOD_TRAINING_0_LOAD19to19;
wire   [20:20]   IOD_TRAINING_0_LOAD20to20;
wire   [21:21]   IOD_TRAINING_0_LOAD21to21;
wire   [22:22]   IOD_TRAINING_0_LOAD22to22;
wire   [23:23]   IOD_TRAINING_0_LOAD23to23;
wire   [24:24]   IOD_TRAINING_0_LOAD24to24;
wire   [25:25]   IOD_TRAINING_0_LOAD25to25;
wire   [26:26]   IOD_TRAINING_0_LOAD26to26;
wire   [27:27]   IOD_TRAINING_0_LOAD27to27;
wire   [28:28]   IOD_TRAINING_0_LOAD28to28;
wire   [29:29]   IOD_TRAINING_0_LOAD29to29;
wire   [30:30]   IOD_TRAINING_0_LOAD30to30;
wire   [31:31]   IOD_TRAINING_0_LOAD31to31;
wire   [32:32]   IOD_TRAINING_0_LOAD32to32;
wire   [33:33]   IOD_TRAINING_0_LOAD33to33;
wire   [34:34]   IOD_TRAINING_0_LOAD34to34;
wire   [35:35]   IOD_TRAINING_0_LOAD35to35;
wire   [0:0]     IOD_TRAINING_0_MOVE0to0;
wire   [1:1]     IOD_TRAINING_0_MOVE1to1;
wire   [2:2]     IOD_TRAINING_0_MOVE2to2;
wire   [3:3]     IOD_TRAINING_0_MOVE3to3;
wire   [4:4]     IOD_TRAINING_0_MOVE4to4;
wire   [5:5]     IOD_TRAINING_0_MOVE5to5;
wire   [6:6]     IOD_TRAINING_0_MOVE6to6;
wire   [7:7]     IOD_TRAINING_0_MOVE7to7;
wire   [8:8]     IOD_TRAINING_0_MOVE8to8;
wire   [9:9]     IOD_TRAINING_0_MOVE9to9;
wire   [10:10]   IOD_TRAINING_0_MOVE10to10;
wire   [11:11]   IOD_TRAINING_0_MOVE11to11;
wire   [12:12]   IOD_TRAINING_0_MOVE12to12;
wire   [13:13]   IOD_TRAINING_0_MOVE13to13;
wire   [14:14]   IOD_TRAINING_0_MOVE14to14;
wire   [15:15]   IOD_TRAINING_0_MOVE15to15;
wire   [16:16]   IOD_TRAINING_0_MOVE16to16;
wire   [17:17]   IOD_TRAINING_0_MOVE17to17;
wire   [18:18]   IOD_TRAINING_0_MOVE18to18;
wire   [19:19]   IOD_TRAINING_0_MOVE19to19;
wire   [20:20]   IOD_TRAINING_0_MOVE20to20;
wire   [21:21]   IOD_TRAINING_0_MOVE21to21;
wire   [22:22]   IOD_TRAINING_0_MOVE22to22;
wire   [23:23]   IOD_TRAINING_0_MOVE23to23;
wire   [24:24]   IOD_TRAINING_0_MOVE24to24;
wire   [25:25]   IOD_TRAINING_0_MOVE25to25;
wire   [26:26]   IOD_TRAINING_0_MOVE26to26;
wire   [27:27]   IOD_TRAINING_0_MOVE27to27;
wire   [28:28]   IOD_TRAINING_0_MOVE28to28;
wire   [29:29]   IOD_TRAINING_0_MOVE29to29;
wire   [30:30]   IOD_TRAINING_0_MOVE30to30;
wire   [31:31]   IOD_TRAINING_0_MOVE31to31;
wire   [32:32]   IOD_TRAINING_0_MOVE32to32;
wire   [33:33]   IOD_TRAINING_0_MOVE33to33;
wire   [34:34]   IOD_TRAINING_0_MOVE34to34;
wire   [35:35]   IOD_TRAINING_0_MOVE35to35;
wire             IOD_TRAINING_0_REFCLK_DELAY_LINE_DIRECTION;
wire             IOD_TRAINING_0_REFCLK_DELAY_LINE_LOAD;
wire             IOD_TRAINING_0_REFCLK_DELAY_LINE_MOVE;
wire             IOD_TRAINING_0_REFCLK_EYE_MONITOR_CLR_FLAGS;
wire   [3:0]     ITER_COUNT_net_0;
wire             LANE_0_CTRL_ARST_N;
wire   [2:0]     LANE_0_CTRL_EYE_MONITOR_WIDTH_OUT;
wire   [2:0]     LANE_0_CTRL_FIFO_RD_PTR;
wire   [2:0]     LANE_0_CTRL_FIFO_WR_PTR;
wire             LANE_0_CTRL_RX_BURST_DETECT;
wire             LANE_0_CTRL_RX_DATA_VALID;
wire             LANE_0_CTRL_RX_DELAY_LINE_OUT_OF_RANGE;
wire   [0:0]     LANE_0_CTRL_RX_DQS_90;
wire             LANE_0_CTRL_RX_SYNC_RST;
wire             LANE_0_CTRL_TX_DELAY_LINE_OUT_OF_RANGE;
wire             LANE_0_CTRL_TX_DQS;
wire             LANE_0_CTRL_TX_DQS_270;
wire             LANE_0_CTRL_TX_SYNC_RST;
wire             LANE_0_IOD_DM_RX_FB;
wire             LANE_0_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_0;
wire             LANE_0_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_1;
wire             LANE_0_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_2;
wire             LANE_0_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_3;
wire             LANE_0_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_4;
wire             LANE_0_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_5;
wire             LANE_0_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_6;
wire             LANE_0_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_7;
wire             LANE_0_IOD_DQ_RX_BYPASS_DATA_0;
wire             LANE_0_IOD_DQ_RX_BYPASS_DATA_1;
wire             LANE_0_IOD_DQ_RX_BYPASS_DATA_2;
wire             LANE_0_IOD_DQ_RX_BYPASS_DATA_3;
wire             LANE_0_IOD_DQ_RX_BYPASS_DATA_4;
wire             LANE_0_IOD_DQ_RX_BYPASS_DATA_5;
wire             LANE_0_IOD_DQ_RX_BYPASS_DATA_6;
wire             LANE_0_IOD_DQ_RX_BYPASS_DATA_7;
wire   [0:0]     LANE_0_IOD_DQ_RX_DATA_00to0;
wire   [1:1]     LANE_0_IOD_DQ_RX_DATA_01to1;
wire   [2:2]     LANE_0_IOD_DQ_RX_DATA_02to2;
wire   [3:3]     LANE_0_IOD_DQ_RX_DATA_03to3;
wire   [4:4]     LANE_0_IOD_DQ_RX_DATA_04to4;
wire   [5:5]     LANE_0_IOD_DQ_RX_DATA_05to5;
wire   [6:6]     LANE_0_IOD_DQ_RX_DATA_06to6;
wire   [7:7]     LANE_0_IOD_DQ_RX_DATA_07to7;
wire   [0:0]     LANE_0_IOD_DQ_RX_DATA_10to0;
wire   [1:1]     LANE_0_IOD_DQ_RX_DATA_11to1;
wire   [2:2]     LANE_0_IOD_DQ_RX_DATA_12to2;
wire   [3:3]     LANE_0_IOD_DQ_RX_DATA_13to3;
wire   [4:4]     LANE_0_IOD_DQ_RX_DATA_14to4;
wire   [5:5]     LANE_0_IOD_DQ_RX_DATA_15to5;
wire   [6:6]     LANE_0_IOD_DQ_RX_DATA_16to6;
wire   [7:7]     LANE_0_IOD_DQ_RX_DATA_17to7;
wire   [0:0]     LANE_0_IOD_DQ_RX_DATA_20to0;
wire   [1:1]     LANE_0_IOD_DQ_RX_DATA_21to1;
wire   [2:2]     LANE_0_IOD_DQ_RX_DATA_22to2;
wire   [3:3]     LANE_0_IOD_DQ_RX_DATA_23to3;
wire   [4:4]     LANE_0_IOD_DQ_RX_DATA_24to4;
wire   [5:5]     LANE_0_IOD_DQ_RX_DATA_25to5;
wire   [6:6]     LANE_0_IOD_DQ_RX_DATA_26to6;
wire   [7:7]     LANE_0_IOD_DQ_RX_DATA_27to7;
wire   [0:0]     LANE_0_IOD_DQ_RX_DATA_30to0;
wire   [1:1]     LANE_0_IOD_DQ_RX_DATA_31to1;
wire   [2:2]     LANE_0_IOD_DQ_RX_DATA_32to2;
wire   [3:3]     LANE_0_IOD_DQ_RX_DATA_33to3;
wire   [4:4]     LANE_0_IOD_DQ_RX_DATA_34to4;
wire   [5:5]     LANE_0_IOD_DQ_RX_DATA_35to5;
wire   [6:6]     LANE_0_IOD_DQ_RX_DATA_36to6;
wire   [7:7]     LANE_0_IOD_DQ_RX_DATA_37to7;
wire   [0:0]     LANE_0_IOD_DQ_RX_DATA_40to0;
wire   [1:1]     LANE_0_IOD_DQ_RX_DATA_41to1;
wire   [2:2]     LANE_0_IOD_DQ_RX_DATA_42to2;
wire   [3:3]     LANE_0_IOD_DQ_RX_DATA_43to3;
wire   [4:4]     LANE_0_IOD_DQ_RX_DATA_44to4;
wire   [5:5]     LANE_0_IOD_DQ_RX_DATA_45to5;
wire   [6:6]     LANE_0_IOD_DQ_RX_DATA_46to6;
wire   [7:7]     LANE_0_IOD_DQ_RX_DATA_47to7;
wire   [0:0]     LANE_0_IOD_DQ_RX_DATA_50to0;
wire   [1:1]     LANE_0_IOD_DQ_RX_DATA_51to1;
wire   [2:2]     LANE_0_IOD_DQ_RX_DATA_52to2;
wire   [3:3]     LANE_0_IOD_DQ_RX_DATA_53to3;
wire   [4:4]     LANE_0_IOD_DQ_RX_DATA_54to4;
wire   [5:5]     LANE_0_IOD_DQ_RX_DATA_55to5;
wire   [6:6]     LANE_0_IOD_DQ_RX_DATA_56to6;
wire   [7:7]     LANE_0_IOD_DQ_RX_DATA_57to7;
wire   [0:0]     LANE_0_IOD_DQ_RX_DATA_60to0;
wire   [1:1]     LANE_0_IOD_DQ_RX_DATA_61to1;
wire   [2:2]     LANE_0_IOD_DQ_RX_DATA_62to2;
wire   [3:3]     LANE_0_IOD_DQ_RX_DATA_63to3;
wire   [4:4]     LANE_0_IOD_DQ_RX_DATA_64to4;
wire   [5:5]     LANE_0_IOD_DQ_RX_DATA_65to5;
wire   [6:6]     LANE_0_IOD_DQ_RX_DATA_66to6;
wire   [7:7]     LANE_0_IOD_DQ_RX_DATA_67to7;
wire   [0:0]     LANE_0_IOD_DQ_RX_DATA_70to0;
wire   [1:1]     LANE_0_IOD_DQ_RX_DATA_71to1;
wire   [2:2]     LANE_0_IOD_DQ_RX_DATA_72to2;
wire   [3:3]     LANE_0_IOD_DQ_RX_DATA_73to3;
wire   [4:4]     LANE_0_IOD_DQ_RX_DATA_74to4;
wire   [5:5]     LANE_0_IOD_DQ_RX_DATA_75to5;
wire   [6:6]     LANE_0_IOD_DQ_RX_DATA_76to6;
wire   [7:7]     LANE_0_IOD_DQ_RX_DATA_77to7;
wire             LANE_0_IOD_DQS_DQS;
wire             LANE_0_IOD_DQS_DQS_N;
wire             LANE_0_IOD_DQSW_TRAINING_DELAY_LINE_OUT_OF_RANGE_0;
wire             LANE_0_IOD_DQSW_TRAINING_EYE_MONITOR_EARLY_0;
wire             LANE_0_IOD_DQSW_TRAINING_EYE_MONITOR_LATE_0;
wire             LANE_0_IOD_DQSW_TRAINING_OE_0;
wire   [0:0]     LANE_0_IOD_DQSW_TRAINING_RX_DATA_00to0;
wire   [1:1]     LANE_0_IOD_DQSW_TRAINING_RX_DATA_01to1;
wire             LANE_0_IOD_DQSW_TRAINING_TX_0;
wire             LANE_0_IOD_READ_TRAINING_DDR_DO_READ;
wire             LANE_0_IOD_READ_TRAINING_DELAY_LINE_OUT_OF_RANGE_0;
wire             LANE_0_IOD_READ_TRAINING_EYE_MONITOR_EARLY_0;
wire             LANE_0_IOD_READ_TRAINING_EYE_MONITOR_LATE_0;
wire   [6:6]     LANE_0_IOD_READ_TRAINING_RX_DATA_06to6;
wire   [7:7]     LANE_0_IOD_READ_TRAINING_RX_DATA_07to7;
wire             LANE_0_IOD_READ_TRAINING_SWITCH;
wire             LANE_1_CTRL_ARST_N;
wire   [2:0]     LANE_1_CTRL_EYE_MONITOR_WIDTH_OUT;
wire   [2:0]     LANE_1_CTRL_FIFO_RD_PTR;
wire   [2:0]     LANE_1_CTRL_FIFO_WR_PTR;
wire             LANE_1_CTRL_RX_BURST_DETECT;
wire             LANE_1_CTRL_RX_DATA_VALID;
wire             LANE_1_CTRL_RX_DELAY_LINE_OUT_OF_RANGE;
wire   [0:0]     LANE_1_CTRL_RX_DQS_90;
wire             LANE_1_CTRL_RX_SYNC_RST;
wire             LANE_1_CTRL_TX_DELAY_LINE_OUT_OF_RANGE;
wire             LANE_1_CTRL_TX_DQS;
wire             LANE_1_CTRL_TX_DQS_270;
wire             LANE_1_CTRL_TX_SYNC_RST;
wire             LANE_1_IOD_DM_RX_FB;
wire             LANE_1_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_0;
wire             LANE_1_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_1;
wire             LANE_1_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_2;
wire             LANE_1_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_3;
wire             LANE_1_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_4;
wire             LANE_1_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_5;
wire             LANE_1_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_6;
wire             LANE_1_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_7;
wire             LANE_1_IOD_DQ_RX_BYPASS_DATA_0;
wire             LANE_1_IOD_DQ_RX_BYPASS_DATA_1;
wire             LANE_1_IOD_DQ_RX_BYPASS_DATA_2;
wire             LANE_1_IOD_DQ_RX_BYPASS_DATA_3;
wire             LANE_1_IOD_DQ_RX_BYPASS_DATA_4;
wire             LANE_1_IOD_DQ_RX_BYPASS_DATA_5;
wire             LANE_1_IOD_DQ_RX_BYPASS_DATA_6;
wire             LANE_1_IOD_DQ_RX_BYPASS_DATA_7;
wire   [0:0]     LANE_1_IOD_DQ_RX_DATA_00to0;
wire   [1:1]     LANE_1_IOD_DQ_RX_DATA_01to1;
wire   [2:2]     LANE_1_IOD_DQ_RX_DATA_02to2;
wire   [3:3]     LANE_1_IOD_DQ_RX_DATA_03to3;
wire   [4:4]     LANE_1_IOD_DQ_RX_DATA_04to4;
wire   [5:5]     LANE_1_IOD_DQ_RX_DATA_05to5;
wire   [6:6]     LANE_1_IOD_DQ_RX_DATA_06to6;
wire   [7:7]     LANE_1_IOD_DQ_RX_DATA_07to7;
wire   [0:0]     LANE_1_IOD_DQ_RX_DATA_10to0;
wire   [1:1]     LANE_1_IOD_DQ_RX_DATA_11to1;
wire   [2:2]     LANE_1_IOD_DQ_RX_DATA_12to2;
wire   [3:3]     LANE_1_IOD_DQ_RX_DATA_13to3;
wire   [4:4]     LANE_1_IOD_DQ_RX_DATA_14to4;
wire   [5:5]     LANE_1_IOD_DQ_RX_DATA_15to5;
wire   [6:6]     LANE_1_IOD_DQ_RX_DATA_16to6;
wire   [7:7]     LANE_1_IOD_DQ_RX_DATA_17to7;
wire   [0:0]     LANE_1_IOD_DQ_RX_DATA_20to0;
wire   [1:1]     LANE_1_IOD_DQ_RX_DATA_21to1;
wire   [2:2]     LANE_1_IOD_DQ_RX_DATA_22to2;
wire   [3:3]     LANE_1_IOD_DQ_RX_DATA_23to3;
wire   [4:4]     LANE_1_IOD_DQ_RX_DATA_24to4;
wire   [5:5]     LANE_1_IOD_DQ_RX_DATA_25to5;
wire   [6:6]     LANE_1_IOD_DQ_RX_DATA_26to6;
wire   [7:7]     LANE_1_IOD_DQ_RX_DATA_27to7;
wire   [0:0]     LANE_1_IOD_DQ_RX_DATA_30to0;
wire   [1:1]     LANE_1_IOD_DQ_RX_DATA_31to1;
wire   [2:2]     LANE_1_IOD_DQ_RX_DATA_32to2;
wire   [3:3]     LANE_1_IOD_DQ_RX_DATA_33to3;
wire   [4:4]     LANE_1_IOD_DQ_RX_DATA_34to4;
wire   [5:5]     LANE_1_IOD_DQ_RX_DATA_35to5;
wire   [6:6]     LANE_1_IOD_DQ_RX_DATA_36to6;
wire   [7:7]     LANE_1_IOD_DQ_RX_DATA_37to7;
wire   [0:0]     LANE_1_IOD_DQ_RX_DATA_40to0;
wire   [1:1]     LANE_1_IOD_DQ_RX_DATA_41to1;
wire   [2:2]     LANE_1_IOD_DQ_RX_DATA_42to2;
wire   [3:3]     LANE_1_IOD_DQ_RX_DATA_43to3;
wire   [4:4]     LANE_1_IOD_DQ_RX_DATA_44to4;
wire   [5:5]     LANE_1_IOD_DQ_RX_DATA_45to5;
wire   [6:6]     LANE_1_IOD_DQ_RX_DATA_46to6;
wire   [7:7]     LANE_1_IOD_DQ_RX_DATA_47to7;
wire   [0:0]     LANE_1_IOD_DQ_RX_DATA_50to0;
wire   [1:1]     LANE_1_IOD_DQ_RX_DATA_51to1;
wire   [2:2]     LANE_1_IOD_DQ_RX_DATA_52to2;
wire   [3:3]     LANE_1_IOD_DQ_RX_DATA_53to3;
wire   [4:4]     LANE_1_IOD_DQ_RX_DATA_54to4;
wire   [5:5]     LANE_1_IOD_DQ_RX_DATA_55to5;
wire   [6:6]     LANE_1_IOD_DQ_RX_DATA_56to6;
wire   [7:7]     LANE_1_IOD_DQ_RX_DATA_57to7;
wire   [0:0]     LANE_1_IOD_DQ_RX_DATA_60to0;
wire   [1:1]     LANE_1_IOD_DQ_RX_DATA_61to1;
wire   [2:2]     LANE_1_IOD_DQ_RX_DATA_62to2;
wire   [3:3]     LANE_1_IOD_DQ_RX_DATA_63to3;
wire   [4:4]     LANE_1_IOD_DQ_RX_DATA_64to4;
wire   [5:5]     LANE_1_IOD_DQ_RX_DATA_65to5;
wire   [6:6]     LANE_1_IOD_DQ_RX_DATA_66to6;
wire   [7:7]     LANE_1_IOD_DQ_RX_DATA_67to7;
wire   [0:0]     LANE_1_IOD_DQ_RX_DATA_70to0;
wire   [1:1]     LANE_1_IOD_DQ_RX_DATA_71to1;
wire   [2:2]     LANE_1_IOD_DQ_RX_DATA_72to2;
wire   [3:3]     LANE_1_IOD_DQ_RX_DATA_73to3;
wire   [4:4]     LANE_1_IOD_DQ_RX_DATA_74to4;
wire   [5:5]     LANE_1_IOD_DQ_RX_DATA_75to5;
wire   [6:6]     LANE_1_IOD_DQ_RX_DATA_76to6;
wire   [7:7]     LANE_1_IOD_DQ_RX_DATA_77to7;
wire             LANE_1_IOD_DQS_DQS;
wire             LANE_1_IOD_DQS_DQS_N;
wire             LANE_1_IOD_DQSW_TRAINING_DELAY_LINE_OUT_OF_RANGE_0;
wire             LANE_1_IOD_DQSW_TRAINING_EYE_MONITOR_EARLY_0;
wire             LANE_1_IOD_DQSW_TRAINING_EYE_MONITOR_LATE_0;
wire             LANE_1_IOD_DQSW_TRAINING_OE_0;
wire   [0:0]     LANE_1_IOD_DQSW_TRAINING_RX_DATA_00to0;
wire   [1:1]     LANE_1_IOD_DQSW_TRAINING_RX_DATA_01to1;
wire             LANE_1_IOD_DQSW_TRAINING_TX_0;
wire             LANE_1_IOD_READ_TRAINING_DDR_DO_READ;
wire             LANE_1_IOD_READ_TRAINING_DELAY_LINE_OUT_OF_RANGE_0;
wire             LANE_1_IOD_READ_TRAINING_EYE_MONITOR_EARLY_0;
wire             LANE_1_IOD_READ_TRAINING_EYE_MONITOR_LATE_0;
wire   [6:6]     LANE_1_IOD_READ_TRAINING_RX_DATA_06to6;
wire   [7:7]     LANE_1_IOD_READ_TRAINING_RX_DATA_07to7;
wire             LANE_1_IOD_READ_TRAINING_SWITCH;
wire             LANE_2_CTRL_ARST_N;
wire   [2:0]     LANE_2_CTRL_EYE_MONITOR_WIDTH_OUT;
wire   [2:0]     LANE_2_CTRL_FIFO_RD_PTR;
wire   [2:0]     LANE_2_CTRL_FIFO_WR_PTR;
wire             LANE_2_CTRL_RX_BURST_DETECT;
wire             LANE_2_CTRL_RX_DATA_VALID;
wire             LANE_2_CTRL_RX_DELAY_LINE_OUT_OF_RANGE;
wire   [0:0]     LANE_2_CTRL_RX_DQS_90;
wire             LANE_2_CTRL_RX_SYNC_RST;
wire             LANE_2_CTRL_TX_DELAY_LINE_OUT_OF_RANGE;
wire             LANE_2_CTRL_TX_DQS;
wire             LANE_2_CTRL_TX_DQS_270;
wire             LANE_2_CTRL_TX_SYNC_RST;
wire             LANE_2_IOD_DM_RX_FB;
wire             LANE_2_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_0;
wire             LANE_2_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_1;
wire             LANE_2_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_2;
wire             LANE_2_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_3;
wire             LANE_2_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_4;
wire             LANE_2_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_5;
wire             LANE_2_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_6;
wire             LANE_2_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_7;
wire             LANE_2_IOD_DQ_RX_BYPASS_DATA_0;
wire             LANE_2_IOD_DQ_RX_BYPASS_DATA_1;
wire             LANE_2_IOD_DQ_RX_BYPASS_DATA_2;
wire             LANE_2_IOD_DQ_RX_BYPASS_DATA_3;
wire             LANE_2_IOD_DQ_RX_BYPASS_DATA_4;
wire             LANE_2_IOD_DQ_RX_BYPASS_DATA_5;
wire             LANE_2_IOD_DQ_RX_BYPASS_DATA_6;
wire             LANE_2_IOD_DQ_RX_BYPASS_DATA_7;
wire   [0:0]     LANE_2_IOD_DQ_RX_DATA_00to0;
wire   [1:1]     LANE_2_IOD_DQ_RX_DATA_01to1;
wire   [2:2]     LANE_2_IOD_DQ_RX_DATA_02to2;
wire   [3:3]     LANE_2_IOD_DQ_RX_DATA_03to3;
wire   [4:4]     LANE_2_IOD_DQ_RX_DATA_04to4;
wire   [5:5]     LANE_2_IOD_DQ_RX_DATA_05to5;
wire   [6:6]     LANE_2_IOD_DQ_RX_DATA_06to6;
wire   [7:7]     LANE_2_IOD_DQ_RX_DATA_07to7;
wire   [0:0]     LANE_2_IOD_DQ_RX_DATA_10to0;
wire   [1:1]     LANE_2_IOD_DQ_RX_DATA_11to1;
wire   [2:2]     LANE_2_IOD_DQ_RX_DATA_12to2;
wire   [3:3]     LANE_2_IOD_DQ_RX_DATA_13to3;
wire   [4:4]     LANE_2_IOD_DQ_RX_DATA_14to4;
wire   [5:5]     LANE_2_IOD_DQ_RX_DATA_15to5;
wire   [6:6]     LANE_2_IOD_DQ_RX_DATA_16to6;
wire   [7:7]     LANE_2_IOD_DQ_RX_DATA_17to7;
wire   [0:0]     LANE_2_IOD_DQ_RX_DATA_20to0;
wire   [1:1]     LANE_2_IOD_DQ_RX_DATA_21to1;
wire   [2:2]     LANE_2_IOD_DQ_RX_DATA_22to2;
wire   [3:3]     LANE_2_IOD_DQ_RX_DATA_23to3;
wire   [4:4]     LANE_2_IOD_DQ_RX_DATA_24to4;
wire   [5:5]     LANE_2_IOD_DQ_RX_DATA_25to5;
wire   [6:6]     LANE_2_IOD_DQ_RX_DATA_26to6;
wire   [7:7]     LANE_2_IOD_DQ_RX_DATA_27to7;
wire   [0:0]     LANE_2_IOD_DQ_RX_DATA_30to0;
wire   [1:1]     LANE_2_IOD_DQ_RX_DATA_31to1;
wire   [2:2]     LANE_2_IOD_DQ_RX_DATA_32to2;
wire   [3:3]     LANE_2_IOD_DQ_RX_DATA_33to3;
wire   [4:4]     LANE_2_IOD_DQ_RX_DATA_34to4;
wire   [5:5]     LANE_2_IOD_DQ_RX_DATA_35to5;
wire   [6:6]     LANE_2_IOD_DQ_RX_DATA_36to6;
wire   [7:7]     LANE_2_IOD_DQ_RX_DATA_37to7;
wire   [0:0]     LANE_2_IOD_DQ_RX_DATA_40to0;
wire   [1:1]     LANE_2_IOD_DQ_RX_DATA_41to1;
wire   [2:2]     LANE_2_IOD_DQ_RX_DATA_42to2;
wire   [3:3]     LANE_2_IOD_DQ_RX_DATA_43to3;
wire   [4:4]     LANE_2_IOD_DQ_RX_DATA_44to4;
wire   [5:5]     LANE_2_IOD_DQ_RX_DATA_45to5;
wire   [6:6]     LANE_2_IOD_DQ_RX_DATA_46to6;
wire   [7:7]     LANE_2_IOD_DQ_RX_DATA_47to7;
wire   [0:0]     LANE_2_IOD_DQ_RX_DATA_50to0;
wire   [1:1]     LANE_2_IOD_DQ_RX_DATA_51to1;
wire   [2:2]     LANE_2_IOD_DQ_RX_DATA_52to2;
wire   [3:3]     LANE_2_IOD_DQ_RX_DATA_53to3;
wire   [4:4]     LANE_2_IOD_DQ_RX_DATA_54to4;
wire   [5:5]     LANE_2_IOD_DQ_RX_DATA_55to5;
wire   [6:6]     LANE_2_IOD_DQ_RX_DATA_56to6;
wire   [7:7]     LANE_2_IOD_DQ_RX_DATA_57to7;
wire   [0:0]     LANE_2_IOD_DQ_RX_DATA_60to0;
wire   [1:1]     LANE_2_IOD_DQ_RX_DATA_61to1;
wire   [2:2]     LANE_2_IOD_DQ_RX_DATA_62to2;
wire   [3:3]     LANE_2_IOD_DQ_RX_DATA_63to3;
wire   [4:4]     LANE_2_IOD_DQ_RX_DATA_64to4;
wire   [5:5]     LANE_2_IOD_DQ_RX_DATA_65to5;
wire   [6:6]     LANE_2_IOD_DQ_RX_DATA_66to6;
wire   [7:7]     LANE_2_IOD_DQ_RX_DATA_67to7;
wire   [0:0]     LANE_2_IOD_DQ_RX_DATA_70to0;
wire   [1:1]     LANE_2_IOD_DQ_RX_DATA_71to1;
wire   [2:2]     LANE_2_IOD_DQ_RX_DATA_72to2;
wire   [3:3]     LANE_2_IOD_DQ_RX_DATA_73to3;
wire   [4:4]     LANE_2_IOD_DQ_RX_DATA_74to4;
wire   [5:5]     LANE_2_IOD_DQ_RX_DATA_75to5;
wire   [6:6]     LANE_2_IOD_DQ_RX_DATA_76to6;
wire   [7:7]     LANE_2_IOD_DQ_RX_DATA_77to7;
wire             LANE_2_IOD_DQS_DQS;
wire             LANE_2_IOD_DQS_DQS_N;
wire             LANE_2_IOD_DQSW_TRAINING_DELAY_LINE_OUT_OF_RANGE_0;
wire             LANE_2_IOD_DQSW_TRAINING_EYE_MONITOR_EARLY_0;
wire             LANE_2_IOD_DQSW_TRAINING_EYE_MONITOR_LATE_0;
wire             LANE_2_IOD_DQSW_TRAINING_OE_0;
wire   [0:0]     LANE_2_IOD_DQSW_TRAINING_RX_DATA_00to0;
wire   [1:1]     LANE_2_IOD_DQSW_TRAINING_RX_DATA_01to1;
wire             LANE_2_IOD_DQSW_TRAINING_TX_0;
wire             LANE_2_IOD_READ_TRAINING_DDR_DO_READ;
wire             LANE_2_IOD_READ_TRAINING_DELAY_LINE_OUT_OF_RANGE_0;
wire             LANE_2_IOD_READ_TRAINING_EYE_MONITOR_EARLY_0;
wire             LANE_2_IOD_READ_TRAINING_EYE_MONITOR_LATE_0;
wire   [6:6]     LANE_2_IOD_READ_TRAINING_RX_DATA_06to6;
wire   [7:7]     LANE_2_IOD_READ_TRAINING_RX_DATA_07to7;
wire             LANE_2_IOD_READ_TRAINING_SWITCH;
wire             LANE_3_CTRL_ARST_N;
wire   [2:0]     LANE_3_CTRL_EYE_MONITOR_WIDTH_OUT;
wire   [2:0]     LANE_3_CTRL_FIFO_RD_PTR;
wire   [2:0]     LANE_3_CTRL_FIFO_WR_PTR;
wire             LANE_3_CTRL_RX_BURST_DETECT;
wire             LANE_3_CTRL_RX_DATA_VALID;
wire             LANE_3_CTRL_RX_DELAY_LINE_OUT_OF_RANGE;
wire   [0:0]     LANE_3_CTRL_RX_DQS_90;
wire             LANE_3_CTRL_RX_SYNC_RST;
wire             LANE_3_CTRL_TX_DELAY_LINE_OUT_OF_RANGE;
wire             LANE_3_CTRL_TX_DQS;
wire             LANE_3_CTRL_TX_DQS_270;
wire             LANE_3_CTRL_TX_SYNC_RST;
wire             LANE_3_IOD_DM_RX_FB;
wire             LANE_3_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_0;
wire             LANE_3_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_1;
wire             LANE_3_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_2;
wire             LANE_3_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_3;
wire             LANE_3_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_4;
wire             LANE_3_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_5;
wire             LANE_3_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_6;
wire             LANE_3_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_7;
wire             LANE_3_IOD_DQ_RX_BYPASS_DATA_0;
wire             LANE_3_IOD_DQ_RX_BYPASS_DATA_1;
wire             LANE_3_IOD_DQ_RX_BYPASS_DATA_2;
wire             LANE_3_IOD_DQ_RX_BYPASS_DATA_3;
wire             LANE_3_IOD_DQ_RX_BYPASS_DATA_4;
wire             LANE_3_IOD_DQ_RX_BYPASS_DATA_5;
wire             LANE_3_IOD_DQ_RX_BYPASS_DATA_6;
wire             LANE_3_IOD_DQ_RX_BYPASS_DATA_7;
wire   [0:0]     LANE_3_IOD_DQ_RX_DATA_00to0;
wire   [1:1]     LANE_3_IOD_DQ_RX_DATA_01to1;
wire   [2:2]     LANE_3_IOD_DQ_RX_DATA_02to2;
wire   [3:3]     LANE_3_IOD_DQ_RX_DATA_03to3;
wire   [4:4]     LANE_3_IOD_DQ_RX_DATA_04to4;
wire   [5:5]     LANE_3_IOD_DQ_RX_DATA_05to5;
wire   [6:6]     LANE_3_IOD_DQ_RX_DATA_06to6;
wire   [7:7]     LANE_3_IOD_DQ_RX_DATA_07to7;
wire   [0:0]     LANE_3_IOD_DQ_RX_DATA_10to0;
wire   [1:1]     LANE_3_IOD_DQ_RX_DATA_11to1;
wire   [2:2]     LANE_3_IOD_DQ_RX_DATA_12to2;
wire   [3:3]     LANE_3_IOD_DQ_RX_DATA_13to3;
wire   [4:4]     LANE_3_IOD_DQ_RX_DATA_14to4;
wire   [5:5]     LANE_3_IOD_DQ_RX_DATA_15to5;
wire   [6:6]     LANE_3_IOD_DQ_RX_DATA_16to6;
wire   [7:7]     LANE_3_IOD_DQ_RX_DATA_17to7;
wire   [0:0]     LANE_3_IOD_DQ_RX_DATA_20to0;
wire   [1:1]     LANE_3_IOD_DQ_RX_DATA_21to1;
wire   [2:2]     LANE_3_IOD_DQ_RX_DATA_22to2;
wire   [3:3]     LANE_3_IOD_DQ_RX_DATA_23to3;
wire   [4:4]     LANE_3_IOD_DQ_RX_DATA_24to4;
wire   [5:5]     LANE_3_IOD_DQ_RX_DATA_25to5;
wire   [6:6]     LANE_3_IOD_DQ_RX_DATA_26to6;
wire   [7:7]     LANE_3_IOD_DQ_RX_DATA_27to7;
wire   [0:0]     LANE_3_IOD_DQ_RX_DATA_30to0;
wire   [1:1]     LANE_3_IOD_DQ_RX_DATA_31to1;
wire   [2:2]     LANE_3_IOD_DQ_RX_DATA_32to2;
wire   [3:3]     LANE_3_IOD_DQ_RX_DATA_33to3;
wire   [4:4]     LANE_3_IOD_DQ_RX_DATA_34to4;
wire   [5:5]     LANE_3_IOD_DQ_RX_DATA_35to5;
wire   [6:6]     LANE_3_IOD_DQ_RX_DATA_36to6;
wire   [7:7]     LANE_3_IOD_DQ_RX_DATA_37to7;
wire   [0:0]     LANE_3_IOD_DQ_RX_DATA_40to0;
wire   [1:1]     LANE_3_IOD_DQ_RX_DATA_41to1;
wire   [2:2]     LANE_3_IOD_DQ_RX_DATA_42to2;
wire   [3:3]     LANE_3_IOD_DQ_RX_DATA_43to3;
wire   [4:4]     LANE_3_IOD_DQ_RX_DATA_44to4;
wire   [5:5]     LANE_3_IOD_DQ_RX_DATA_45to5;
wire   [6:6]     LANE_3_IOD_DQ_RX_DATA_46to6;
wire   [7:7]     LANE_3_IOD_DQ_RX_DATA_47to7;
wire   [0:0]     LANE_3_IOD_DQ_RX_DATA_50to0;
wire   [1:1]     LANE_3_IOD_DQ_RX_DATA_51to1;
wire   [2:2]     LANE_3_IOD_DQ_RX_DATA_52to2;
wire   [3:3]     LANE_3_IOD_DQ_RX_DATA_53to3;
wire   [4:4]     LANE_3_IOD_DQ_RX_DATA_54to4;
wire   [5:5]     LANE_3_IOD_DQ_RX_DATA_55to5;
wire   [6:6]     LANE_3_IOD_DQ_RX_DATA_56to6;
wire   [7:7]     LANE_3_IOD_DQ_RX_DATA_57to7;
wire   [0:0]     LANE_3_IOD_DQ_RX_DATA_60to0;
wire   [1:1]     LANE_3_IOD_DQ_RX_DATA_61to1;
wire   [2:2]     LANE_3_IOD_DQ_RX_DATA_62to2;
wire   [3:3]     LANE_3_IOD_DQ_RX_DATA_63to3;
wire   [4:4]     LANE_3_IOD_DQ_RX_DATA_64to4;
wire   [5:5]     LANE_3_IOD_DQ_RX_DATA_65to5;
wire   [6:6]     LANE_3_IOD_DQ_RX_DATA_66to6;
wire   [7:7]     LANE_3_IOD_DQ_RX_DATA_67to7;
wire   [0:0]     LANE_3_IOD_DQ_RX_DATA_70to0;
wire   [1:1]     LANE_3_IOD_DQ_RX_DATA_71to1;
wire   [2:2]     LANE_3_IOD_DQ_RX_DATA_72to2;
wire   [3:3]     LANE_3_IOD_DQ_RX_DATA_73to3;
wire   [4:4]     LANE_3_IOD_DQ_RX_DATA_74to4;
wire   [5:5]     LANE_3_IOD_DQ_RX_DATA_75to5;
wire   [6:6]     LANE_3_IOD_DQ_RX_DATA_76to6;
wire   [7:7]     LANE_3_IOD_DQ_RX_DATA_77to7;
wire             LANE_3_IOD_DQS_DQS;
wire             LANE_3_IOD_DQS_DQS_N;
wire             LANE_3_IOD_DQSW_TRAINING_DELAY_LINE_OUT_OF_RANGE_0;
wire             LANE_3_IOD_DQSW_TRAINING_EYE_MONITOR_EARLY_0;
wire             LANE_3_IOD_DQSW_TRAINING_EYE_MONITOR_LATE_0;
wire             LANE_3_IOD_DQSW_TRAINING_OE_0;
wire   [0:0]     LANE_3_IOD_DQSW_TRAINING_RX_DATA_00to0;
wire   [1:1]     LANE_3_IOD_DQSW_TRAINING_RX_DATA_01to1;
wire             LANE_3_IOD_DQSW_TRAINING_TX_0;
wire             LANE_3_IOD_READ_TRAINING_DDR_DO_READ;
wire             LANE_3_IOD_READ_TRAINING_DELAY_LINE_OUT_OF_RANGE_0;
wire             LANE_3_IOD_READ_TRAINING_EYE_MONITOR_EARLY_0;
wire             LANE_3_IOD_READ_TRAINING_EYE_MONITOR_LATE_0;
wire   [6:6]     LANE_3_IOD_READ_TRAINING_RX_DATA_06to6;
wire   [7:7]     LANE_3_IOD_READ_TRAINING_RX_DATA_07to7;
wire             LANE_3_IOD_READ_TRAINING_SWITCH;
wire             LANECTRL_ADDR_CMD_0_ARST_N;
wire             LANECTRL_ADDR_CMD_0_RX_SYNC_RST;
wire             LANECTRL_ADDR_CMD_0_TX_DQS_270;
wire             LANECTRL_ADDR_CMD_0_TX_SYNC_RST;
wire   [0:0]     LOADPHS_B_net_0;
wire             OB_A_12_Y;
wire             OB_DIFF_CK0_Y;
wire   [0:0]     ODT_net_0;
wire             PCLK;
wire             PLL_LOCK;
wire   [0:0]     RAS_N_net_0;
wire   [9:0]     RDGATE_MIN_READS_THRESHOLD;
wire             REF_CLK;
wire   [0:0]     RESET_N_net_0;
wire             SHIELD0_net_0;
wire             SHIELD1_net_0;
wire             SHIELD2_net_0;
wire             SHIELD3_net_0;
wire             SKIP_BCLK_TRN;
wire             SKIP_CA_TRN;
wire             SKIP_DQSW_TRN;
wire             SKIP_RDLVL_TRN;
wire             SKIP_VREF_TRAINING;
wire             SKIP_WRLVL_TRN;
wire             SYNC_SYS_RST_N_net_0;
wire             SYS_CLK;
wire             SYS_RST_N;
wire   [0:0]     VCO_PHSEL_BCLK90_SEL_net_0;
wire   [0:0]     VCO_PHSEL_BCLK_SEL_net_0;
wire             VCO_PHSEL_REFCLK_SEL_net_0;
wire   [0:0]     VCO_PHSEL_ROTATE_net_0;
wire   [6:0]     VREF_MR6_VALUE;
wire   [0:0]     WE_N_net_0;
wire   [7:0]     WRCAL_WRITE_COUNTER_VALUE;
wire   [6:0]     WRLVL_TAP_OFFSET;
wire             CODE_UPDATE_net_1;
wire   [0:0]     LOADPHS_B_net_1;
wire   [0:0]     VCO_PHSEL_BCLK_SEL_net_1;
wire   [0:0]     VCO_PHSEL_BCLK90_SEL_net_1;
wire             VCO_PHSEL_REFCLK_SEL_net_1;
wire   [0:0]     VCO_PHSEL_ROTATE_net_1;
wire   [63:0]    DFI_RDDATA_W0_net_1;
wire   [0:0]     DFI_RDDATA_VALID_W0_net_1;
wire   [1:1]     DFI_RDDATA_VALID_W0_net_2;
wire   [2:2]     DFI_RDDATA_VALID_W0_net_3;
wire   [3:3]     DFI_RDDATA_VALID_W0_net_4;
wire   [63:0]    DFI_RDDATA_W1_net_1;
wire   [0:0]     DFI_RDDATA_VALID_W1_net_1;
wire   [1:1]     DFI_RDDATA_VALID_W1_net_2;
wire   [2:2]     DFI_RDDATA_VALID_W1_net_3;
wire   [3:3]     DFI_RDDATA_VALID_W1_net_4;
wire   [63:0]    DFI_RDDATA_W2_net_1;
wire   [0:0]     DFI_RDDATA_VALID_W2_net_1;
wire   [1:1]     DFI_RDDATA_VALID_W2_net_2;
wire   [2:2]     DFI_RDDATA_VALID_W2_net_3;
wire   [3:3]     DFI_RDDATA_VALID_W2_net_4;
wire   [63:0]    DFI_RDDATA_W3_net_1;
wire   [0:0]     DFI_RDDATA_VALID_W3_net_1;
wire   [1:1]     DFI_RDDATA_VALID_W3_net_2;
wire   [2:2]     DFI_RDDATA_VALID_W3_net_3;
wire   [3:3]     DFI_RDDATA_VALID_W3_net_4;
wire   [3:0]     DFI_RDLVL_RESP_net_1;
wire   [3:0]     DFI_WRLVL_RESP_net_1;
wire             DFI_INIT_COMPLETE_net_1;
wire             DFI_TRAINING_COMPLETE_net_1;
wire   [0:0]     DM_N_net_1;
wire   [1:1]     DM_N_0_net_0;
wire   [2:2]     DM_N_1_net_0;
wire   [3:3]     DM_N_2_net_0;
wire             CKE_net_1;
wire             CS_N_net_1;
wire             ODT_net_1;
wire             RAS_N_net_1;
wire             CAS_N_net_1;
wire             WE_N_net_1;
wire             ACT_N_net_1;
wire   [1:0]     BG_net_1;
wire   [1:0]     BA_net_1;
wire             RESET_N_net_1;
wire   [0:0]     A_net_1;
wire   [10:10]   A_9_net_0;
wire   [11:11]   A_10_net_0;
wire   [12:12]   A_11_net_0;
wire   [13:13]   A_12_net_0;
wire   [1:1]     A_0_net_0;
wire   [2:2]     A_1_net_0;
wire   [3:3]     A_2_net_0;
wire   [4:4]     A_3_net_0;
wire   [5:5]     A_4_net_0;
wire   [6:6]     A_5_net_0;
wire   [7:7]     A_6_net_0;
wire   [8:8]     A_7_net_0;
wire   [9:9]     A_8_net_0;
wire             CK0_net_1;
wire             CK0_N_net_1;
wire             SHIELD0_net_1;
wire             SHIELD1_net_1;
wire             SHIELD2_net_1;
wire             SHIELD3_net_1;
wire   [7:0]     APB_DEBUG_PRDATA_net_0;
wire             APB_DEBUG_PREADY_net_0;
wire             CAL_INIT_MR_W_REQ_net_1;
wire   [7:0]     CAL_INIT_MR_ADDR_net_1;
wire   [17:0]    CAL_INIT_MR_WR_DATA_net_1;
wire   [17:0]    CAL_INIT_MR_WR_MASK_net_1;
wire   [1:0]     CAL_INIT_CS_net_1;
wire             CTRLR_READY_OUT_net_1;
wire   [3:0]     ITER_COUNT_net_1;
wire             CAL_L_R_REQ_net_1;
wire             CAL_L_W_REQ_net_1;
wire   [255:0]   CAL_L_DATAIN_net_1;
wire   [31:0]    CAL_L_DM_IN_net_1;
wire             CAL_SELECT_net_1;
wire   [0:0]     DFI_RDDATA_W0_slice_0;
wire   [10:10]   DFI_RDDATA_W0_slice_1;
wire   [11:11]   DFI_RDDATA_W0_slice_2;
wire   [12:12]   DFI_RDDATA_W0_slice_3;
wire   [13:13]   DFI_RDDATA_W0_slice_4;
wire   [14:14]   DFI_RDDATA_W0_slice_5;
wire   [15:15]   DFI_RDDATA_W0_slice_6;
wire   [16:16]   DFI_RDDATA_W0_slice_7;
wire   [17:17]   DFI_RDDATA_W0_slice_8;
wire   [18:18]   DFI_RDDATA_W0_slice_9;
wire   [19:19]   DFI_RDDATA_W0_slice_10;
wire   [1:1]     DFI_RDDATA_W0_slice_11;
wire   [20:20]   DFI_RDDATA_W0_slice_12;
wire   [21:21]   DFI_RDDATA_W0_slice_13;
wire   [22:22]   DFI_RDDATA_W0_slice_14;
wire   [23:23]   DFI_RDDATA_W0_slice_15;
wire   [24:24]   DFI_RDDATA_W0_slice_16;
wire   [25:25]   DFI_RDDATA_W0_slice_17;
wire   [26:26]   DFI_RDDATA_W0_slice_18;
wire   [27:27]   DFI_RDDATA_W0_slice_19;
wire   [28:28]   DFI_RDDATA_W0_slice_20;
wire   [29:29]   DFI_RDDATA_W0_slice_21;
wire   [2:2]     DFI_RDDATA_W0_slice_22;
wire   [30:30]   DFI_RDDATA_W0_slice_23;
wire   [31:31]   DFI_RDDATA_W0_slice_24;
wire   [32:32]   DFI_RDDATA_W0_slice_25;
wire   [33:33]   DFI_RDDATA_W0_slice_26;
wire   [34:34]   DFI_RDDATA_W0_slice_27;
wire   [35:35]   DFI_RDDATA_W0_slice_28;
wire   [36:36]   DFI_RDDATA_W0_slice_29;
wire   [37:37]   DFI_RDDATA_W0_slice_30;
wire   [38:38]   DFI_RDDATA_W0_slice_31;
wire   [39:39]   DFI_RDDATA_W0_slice_32;
wire   [3:3]     DFI_RDDATA_W0_slice_33;
wire   [40:40]   DFI_RDDATA_W0_slice_34;
wire   [41:41]   DFI_RDDATA_W0_slice_35;
wire   [42:42]   DFI_RDDATA_W0_slice_36;
wire   [43:43]   DFI_RDDATA_W0_slice_37;
wire   [44:44]   DFI_RDDATA_W0_slice_38;
wire   [45:45]   DFI_RDDATA_W0_slice_39;
wire   [46:46]   DFI_RDDATA_W0_slice_40;
wire   [47:47]   DFI_RDDATA_W0_slice_41;
wire   [48:48]   DFI_RDDATA_W0_slice_42;
wire   [49:49]   DFI_RDDATA_W0_slice_43;
wire   [4:4]     DFI_RDDATA_W0_slice_44;
wire   [50:50]   DFI_RDDATA_W0_slice_45;
wire   [51:51]   DFI_RDDATA_W0_slice_46;
wire   [52:52]   DFI_RDDATA_W0_slice_47;
wire   [53:53]   DFI_RDDATA_W0_slice_48;
wire   [54:54]   DFI_RDDATA_W0_slice_49;
wire   [55:55]   DFI_RDDATA_W0_slice_50;
wire   [56:56]   DFI_RDDATA_W0_slice_51;
wire   [57:57]   DFI_RDDATA_W0_slice_52;
wire   [58:58]   DFI_RDDATA_W0_slice_53;
wire   [59:59]   DFI_RDDATA_W0_slice_54;
wire   [5:5]     DFI_RDDATA_W0_slice_55;
wire   [60:60]   DFI_RDDATA_W0_slice_56;
wire   [61:61]   DFI_RDDATA_W0_slice_57;
wire   [62:62]   DFI_RDDATA_W0_slice_58;
wire   [63:63]   DFI_RDDATA_W0_slice_59;
wire   [6:6]     DFI_RDDATA_W0_slice_60;
wire   [7:7]     DFI_RDDATA_W0_slice_61;
wire   [8:8]     DFI_RDDATA_W0_slice_62;
wire   [9:9]     DFI_RDDATA_W0_slice_63;
wire   [0:0]     DFI_RDDATA_W1_slice_0;
wire   [10:10]   DFI_RDDATA_W1_slice_1;
wire   [11:11]   DFI_RDDATA_W1_slice_2;
wire   [12:12]   DFI_RDDATA_W1_slice_3;
wire   [13:13]   DFI_RDDATA_W1_slice_4;
wire   [14:14]   DFI_RDDATA_W1_slice_5;
wire   [15:15]   DFI_RDDATA_W1_slice_6;
wire   [16:16]   DFI_RDDATA_W1_slice_7;
wire   [17:17]   DFI_RDDATA_W1_slice_8;
wire   [18:18]   DFI_RDDATA_W1_slice_9;
wire   [19:19]   DFI_RDDATA_W1_slice_10;
wire   [1:1]     DFI_RDDATA_W1_slice_11;
wire   [20:20]   DFI_RDDATA_W1_slice_12;
wire   [21:21]   DFI_RDDATA_W1_slice_13;
wire   [22:22]   DFI_RDDATA_W1_slice_14;
wire   [23:23]   DFI_RDDATA_W1_slice_15;
wire   [24:24]   DFI_RDDATA_W1_slice_16;
wire   [25:25]   DFI_RDDATA_W1_slice_17;
wire   [26:26]   DFI_RDDATA_W1_slice_18;
wire   [27:27]   DFI_RDDATA_W1_slice_19;
wire   [28:28]   DFI_RDDATA_W1_slice_20;
wire   [29:29]   DFI_RDDATA_W1_slice_21;
wire   [2:2]     DFI_RDDATA_W1_slice_22;
wire   [30:30]   DFI_RDDATA_W1_slice_23;
wire   [31:31]   DFI_RDDATA_W1_slice_24;
wire   [32:32]   DFI_RDDATA_W1_slice_25;
wire   [33:33]   DFI_RDDATA_W1_slice_26;
wire   [34:34]   DFI_RDDATA_W1_slice_27;
wire   [35:35]   DFI_RDDATA_W1_slice_28;
wire   [36:36]   DFI_RDDATA_W1_slice_29;
wire   [37:37]   DFI_RDDATA_W1_slice_30;
wire   [38:38]   DFI_RDDATA_W1_slice_31;
wire   [39:39]   DFI_RDDATA_W1_slice_32;
wire   [3:3]     DFI_RDDATA_W1_slice_33;
wire   [40:40]   DFI_RDDATA_W1_slice_34;
wire   [41:41]   DFI_RDDATA_W1_slice_35;
wire   [42:42]   DFI_RDDATA_W1_slice_36;
wire   [43:43]   DFI_RDDATA_W1_slice_37;
wire   [44:44]   DFI_RDDATA_W1_slice_38;
wire   [45:45]   DFI_RDDATA_W1_slice_39;
wire   [46:46]   DFI_RDDATA_W1_slice_40;
wire   [47:47]   DFI_RDDATA_W1_slice_41;
wire   [48:48]   DFI_RDDATA_W1_slice_42;
wire   [49:49]   DFI_RDDATA_W1_slice_43;
wire   [4:4]     DFI_RDDATA_W1_slice_44;
wire   [50:50]   DFI_RDDATA_W1_slice_45;
wire   [51:51]   DFI_RDDATA_W1_slice_46;
wire   [52:52]   DFI_RDDATA_W1_slice_47;
wire   [53:53]   DFI_RDDATA_W1_slice_48;
wire   [54:54]   DFI_RDDATA_W1_slice_49;
wire   [55:55]   DFI_RDDATA_W1_slice_50;
wire   [56:56]   DFI_RDDATA_W1_slice_51;
wire   [57:57]   DFI_RDDATA_W1_slice_52;
wire   [58:58]   DFI_RDDATA_W1_slice_53;
wire   [59:59]   DFI_RDDATA_W1_slice_54;
wire   [5:5]     DFI_RDDATA_W1_slice_55;
wire   [60:60]   DFI_RDDATA_W1_slice_56;
wire   [61:61]   DFI_RDDATA_W1_slice_57;
wire   [62:62]   DFI_RDDATA_W1_slice_58;
wire   [63:63]   DFI_RDDATA_W1_slice_59;
wire   [6:6]     DFI_RDDATA_W1_slice_60;
wire   [7:7]     DFI_RDDATA_W1_slice_61;
wire   [8:8]     DFI_RDDATA_W1_slice_62;
wire   [9:9]     DFI_RDDATA_W1_slice_63;
wire   [0:0]     DFI_RDDATA_W2_slice_0;
wire   [10:10]   DFI_RDDATA_W2_slice_1;
wire   [11:11]   DFI_RDDATA_W2_slice_2;
wire   [12:12]   DFI_RDDATA_W2_slice_3;
wire   [13:13]   DFI_RDDATA_W2_slice_4;
wire   [14:14]   DFI_RDDATA_W2_slice_5;
wire   [15:15]   DFI_RDDATA_W2_slice_6;
wire   [16:16]   DFI_RDDATA_W2_slice_7;
wire   [17:17]   DFI_RDDATA_W2_slice_8;
wire   [18:18]   DFI_RDDATA_W2_slice_9;
wire   [19:19]   DFI_RDDATA_W2_slice_10;
wire   [1:1]     DFI_RDDATA_W2_slice_11;
wire   [20:20]   DFI_RDDATA_W2_slice_12;
wire   [21:21]   DFI_RDDATA_W2_slice_13;
wire   [22:22]   DFI_RDDATA_W2_slice_14;
wire   [23:23]   DFI_RDDATA_W2_slice_15;
wire   [24:24]   DFI_RDDATA_W2_slice_16;
wire   [25:25]   DFI_RDDATA_W2_slice_17;
wire   [26:26]   DFI_RDDATA_W2_slice_18;
wire   [27:27]   DFI_RDDATA_W2_slice_19;
wire   [28:28]   DFI_RDDATA_W2_slice_20;
wire   [29:29]   DFI_RDDATA_W2_slice_21;
wire   [2:2]     DFI_RDDATA_W2_slice_22;
wire   [30:30]   DFI_RDDATA_W2_slice_23;
wire   [31:31]   DFI_RDDATA_W2_slice_24;
wire   [32:32]   DFI_RDDATA_W2_slice_25;
wire   [33:33]   DFI_RDDATA_W2_slice_26;
wire   [34:34]   DFI_RDDATA_W2_slice_27;
wire   [35:35]   DFI_RDDATA_W2_slice_28;
wire   [36:36]   DFI_RDDATA_W2_slice_29;
wire   [37:37]   DFI_RDDATA_W2_slice_30;
wire   [38:38]   DFI_RDDATA_W2_slice_31;
wire   [39:39]   DFI_RDDATA_W2_slice_32;
wire   [3:3]     DFI_RDDATA_W2_slice_33;
wire   [40:40]   DFI_RDDATA_W2_slice_34;
wire   [41:41]   DFI_RDDATA_W2_slice_35;
wire   [42:42]   DFI_RDDATA_W2_slice_36;
wire   [43:43]   DFI_RDDATA_W2_slice_37;
wire   [44:44]   DFI_RDDATA_W2_slice_38;
wire   [45:45]   DFI_RDDATA_W2_slice_39;
wire   [46:46]   DFI_RDDATA_W2_slice_40;
wire   [47:47]   DFI_RDDATA_W2_slice_41;
wire   [48:48]   DFI_RDDATA_W2_slice_42;
wire   [49:49]   DFI_RDDATA_W2_slice_43;
wire   [4:4]     DFI_RDDATA_W2_slice_44;
wire   [50:50]   DFI_RDDATA_W2_slice_45;
wire   [51:51]   DFI_RDDATA_W2_slice_46;
wire   [52:52]   DFI_RDDATA_W2_slice_47;
wire   [53:53]   DFI_RDDATA_W2_slice_48;
wire   [54:54]   DFI_RDDATA_W2_slice_49;
wire   [55:55]   DFI_RDDATA_W2_slice_50;
wire   [56:56]   DFI_RDDATA_W2_slice_51;
wire   [57:57]   DFI_RDDATA_W2_slice_52;
wire   [58:58]   DFI_RDDATA_W2_slice_53;
wire   [59:59]   DFI_RDDATA_W2_slice_54;
wire   [5:5]     DFI_RDDATA_W2_slice_55;
wire   [60:60]   DFI_RDDATA_W2_slice_56;
wire   [61:61]   DFI_RDDATA_W2_slice_57;
wire   [62:62]   DFI_RDDATA_W2_slice_58;
wire   [63:63]   DFI_RDDATA_W2_slice_59;
wire   [6:6]     DFI_RDDATA_W2_slice_60;
wire   [7:7]     DFI_RDDATA_W2_slice_61;
wire   [8:8]     DFI_RDDATA_W2_slice_62;
wire   [9:9]     DFI_RDDATA_W2_slice_63;
wire   [0:0]     DFI_RDDATA_W3_slice_0;
wire   [10:10]   DFI_RDDATA_W3_slice_1;
wire   [11:11]   DFI_RDDATA_W3_slice_2;
wire   [12:12]   DFI_RDDATA_W3_slice_3;
wire   [13:13]   DFI_RDDATA_W3_slice_4;
wire   [14:14]   DFI_RDDATA_W3_slice_5;
wire   [15:15]   DFI_RDDATA_W3_slice_6;
wire   [16:16]   DFI_RDDATA_W3_slice_7;
wire   [17:17]   DFI_RDDATA_W3_slice_8;
wire   [18:18]   DFI_RDDATA_W3_slice_9;
wire   [19:19]   DFI_RDDATA_W3_slice_10;
wire   [1:1]     DFI_RDDATA_W3_slice_11;
wire   [20:20]   DFI_RDDATA_W3_slice_12;
wire   [21:21]   DFI_RDDATA_W3_slice_13;
wire   [22:22]   DFI_RDDATA_W3_slice_14;
wire   [23:23]   DFI_RDDATA_W3_slice_15;
wire   [24:24]   DFI_RDDATA_W3_slice_16;
wire   [25:25]   DFI_RDDATA_W3_slice_17;
wire   [26:26]   DFI_RDDATA_W3_slice_18;
wire   [27:27]   DFI_RDDATA_W3_slice_19;
wire   [28:28]   DFI_RDDATA_W3_slice_20;
wire   [29:29]   DFI_RDDATA_W3_slice_21;
wire   [2:2]     DFI_RDDATA_W3_slice_22;
wire   [30:30]   DFI_RDDATA_W3_slice_23;
wire   [31:31]   DFI_RDDATA_W3_slice_24;
wire   [32:32]   DFI_RDDATA_W3_slice_25;
wire   [33:33]   DFI_RDDATA_W3_slice_26;
wire   [34:34]   DFI_RDDATA_W3_slice_27;
wire   [35:35]   DFI_RDDATA_W3_slice_28;
wire   [36:36]   DFI_RDDATA_W3_slice_29;
wire   [37:37]   DFI_RDDATA_W3_slice_30;
wire   [38:38]   DFI_RDDATA_W3_slice_31;
wire   [39:39]   DFI_RDDATA_W3_slice_32;
wire   [3:3]     DFI_RDDATA_W3_slice_33;
wire   [40:40]   DFI_RDDATA_W3_slice_34;
wire   [41:41]   DFI_RDDATA_W3_slice_35;
wire   [42:42]   DFI_RDDATA_W3_slice_36;
wire   [43:43]   DFI_RDDATA_W3_slice_37;
wire   [44:44]   DFI_RDDATA_W3_slice_38;
wire   [45:45]   DFI_RDDATA_W3_slice_39;
wire   [46:46]   DFI_RDDATA_W3_slice_40;
wire   [47:47]   DFI_RDDATA_W3_slice_41;
wire   [48:48]   DFI_RDDATA_W3_slice_42;
wire   [49:49]   DFI_RDDATA_W3_slice_43;
wire   [4:4]     DFI_RDDATA_W3_slice_44;
wire   [50:50]   DFI_RDDATA_W3_slice_45;
wire   [51:51]   DFI_RDDATA_W3_slice_46;
wire   [52:52]   DFI_RDDATA_W3_slice_47;
wire   [53:53]   DFI_RDDATA_W3_slice_48;
wire   [54:54]   DFI_RDDATA_W3_slice_49;
wire   [55:55]   DFI_RDDATA_W3_slice_50;
wire   [56:56]   DFI_RDDATA_W3_slice_51;
wire   [57:57]   DFI_RDDATA_W3_slice_52;
wire   [58:58]   DFI_RDDATA_W3_slice_53;
wire   [59:59]   DFI_RDDATA_W3_slice_54;
wire   [5:5]     DFI_RDDATA_W3_slice_55;
wire   [60:60]   DFI_RDDATA_W3_slice_56;
wire   [61:61]   DFI_RDDATA_W3_slice_57;
wire   [62:62]   DFI_RDDATA_W3_slice_58;
wire   [63:63]   DFI_RDDATA_W3_slice_59;
wire   [6:6]     DFI_RDDATA_W3_slice_60;
wire   [7:7]     DFI_RDDATA_W3_slice_61;
wire   [8:8]     DFI_RDDATA_W3_slice_62;
wire   [9:9]     DFI_RDDATA_W3_slice_63;
wire   [0:0]     DFI_WRLVL_RESP_slice_0;
wire   [1:1]     DFI_WRLVL_RESP_slice_1;
wire   [2:2]     DFI_WRLVL_RESP_slice_2;
wire   [3:3]     DFI_WRLVL_RESP_slice_3;
wire   [0:0]     RX_DATA_0_slice_0;
wire   [1:1]     RX_DATA_0_slice_1;
wire   [2:2]     RX_DATA_0_slice_2;
wire   [1:1]     RX_DATA_0_slice_3;
wire   [3:3]     RX_DATA_0_slice_4;
wire   [5:5]     RX_DATA_0_slice_5;
wire   [7:7]     RX_DATA_0_slice_6;
wire   [0:0]     RX_DATA_0_slice_7;
wire   [1:1]     RX_DATA_0_slice_8;
wire   [2:2]     RX_DATA_0_slice_9;
wire   [3:3]     RX_DATA_0_slice_10;
wire   [4:4]     RX_DATA_0_slice_11;
wire   [5:5]     RX_DATA_0_slice_12;
wire   [7:7]     RX_DATA_0_slice_13;
wire   [0:0]     ODT_DYN_LANE_slice_0;
wire   [1:1]     ODT_DYN_LANE_slice_1;
wire   [2:2]     ODT_DYN_LANE_slice_2;
wire   [3:3]     ODT_DYN_LANE_slice_3;
wire   [0:0]     IOG_WRDATA_MASK_P0_slice_0;
wire   [1:1]     IOG_WRDATA_MASK_P0_slice_1;
wire   [2:2]     IOG_WRDATA_MASK_P0_slice_2;
wire   [3:3]     IOG_WRDATA_MASK_P0_slice_3;
wire   [4:4]     IOG_WRDATA_MASK_P0_slice_4;
wire   [5:5]     IOG_WRDATA_MASK_P0_slice_5;
wire   [6:6]     IOG_WRDATA_MASK_P0_slice_6;
wire   [7:7]     IOG_WRDATA_MASK_P0_slice_7;
wire   [0:0]     IOG_WRDATA_MASK_P1_slice_0;
wire   [1:1]     IOG_WRDATA_MASK_P1_slice_1;
wire   [2:2]     IOG_WRDATA_MASK_P1_slice_2;
wire   [3:3]     IOG_WRDATA_MASK_P1_slice_3;
wire   [4:4]     IOG_WRDATA_MASK_P1_slice_4;
wire   [5:5]     IOG_WRDATA_MASK_P1_slice_5;
wire   [6:6]     IOG_WRDATA_MASK_P1_slice_6;
wire   [7:7]     IOG_WRDATA_MASK_P1_slice_7;
wire   [0:0]     IOG_WRDATA_MASK_P2_slice_0;
wire   [1:1]     IOG_WRDATA_MASK_P2_slice_1;
wire   [2:2]     IOG_WRDATA_MASK_P2_slice_2;
wire   [3:3]     IOG_WRDATA_MASK_P2_slice_3;
wire   [4:4]     IOG_WRDATA_MASK_P2_slice_4;
wire   [5:5]     IOG_WRDATA_MASK_P2_slice_5;
wire   [6:6]     IOG_WRDATA_MASK_P2_slice_6;
wire   [7:7]     IOG_WRDATA_MASK_P2_slice_7;
wire   [0:0]     IOG_WRDATA_MASK_P3_slice_0;
wire   [1:1]     IOG_WRDATA_MASK_P3_slice_1;
wire   [2:2]     IOG_WRDATA_MASK_P3_slice_2;
wire   [3:3]     IOG_WRDATA_MASK_P3_slice_3;
wire   [4:4]     IOG_WRDATA_MASK_P3_slice_4;
wire   [5:5]     IOG_WRDATA_MASK_P3_slice_5;
wire   [6:6]     IOG_WRDATA_MASK_P3_slice_6;
wire   [7:7]     IOG_WRDATA_MASK_P3_slice_7;
wire   [14:14]   IOG_ADDRESS_P0_slice_0;
wire   [15:15]   IOG_ADDRESS_P0_slice_1;
wire   [16:16]   IOG_ADDRESS_P0_slice_2;
wire   [17:17]   IOG_ADDRESS_P0_slice_3;
wire   [18:18]   IOG_ADDRESS_P0_slice_4;
wire   [19:19]   IOG_ADDRESS_P0_slice_5;
wire   [14:14]   IOG_ADDRESS_P1_slice_0;
wire   [15:15]   IOG_ADDRESS_P1_slice_1;
wire   [16:16]   IOG_ADDRESS_P1_slice_2;
wire   [17:17]   IOG_ADDRESS_P1_slice_3;
wire   [18:18]   IOG_ADDRESS_P1_slice_4;
wire   [19:19]   IOG_ADDRESS_P1_slice_5;
wire   [14:14]   IOG_ADDRESS_P2_slice_0;
wire   [15:15]   IOG_ADDRESS_P2_slice_1;
wire   [16:16]   IOG_ADDRESS_P2_slice_2;
wire   [17:17]   IOG_ADDRESS_P2_slice_3;
wire   [18:18]   IOG_ADDRESS_P2_slice_4;
wire   [19:19]   IOG_ADDRESS_P2_slice_5;
wire   [14:14]   IOG_ADDRESS_P3_slice_0;
wire   [15:15]   IOG_ADDRESS_P3_slice_1;
wire   [16:16]   IOG_ADDRESS_P3_slice_2;
wire   [17:17]   IOG_ADDRESS_P3_slice_3;
wire   [18:18]   IOG_ADDRESS_P3_slice_4;
wire   [19:19]   IOG_ADDRESS_P3_slice_5;
wire   [2:2]     DFI_BANK_P0_OUT_slice_0;
wire   [2:2]     DFI_BANK_P1_OUT_slice_0;
wire   [2:2]     DFI_BANK_P2_OUT_slice_0;
wire   [2:2]     DFI_BANK_P3_OUT_slice_0;
wire   [0:0]     RX_DATA_0_slice_14;
wire   [1:1]     RX_DATA_0_slice_15;
wire   [2:2]     RX_DATA_0_slice_16;
wire   [3:3]     RX_DATA_0_slice_17;
wire   [4:4]     RX_DATA_0_slice_18;
wire   [5:5]     RX_DATA_0_slice_19;
wire   [0:0]     RX_DATA_0_slice_20;
wire   [1:1]     RX_DATA_0_slice_21;
wire   [2:2]     RX_DATA_0_slice_22;
wire   [3:3]     RX_DATA_0_slice_23;
wire   [4:4]     RX_DATA_0_slice_24;
wire   [5:5]     RX_DATA_0_slice_25;
wire   [0:0]     RX_DATA_0_slice_26;
wire   [1:1]     RX_DATA_0_slice_27;
wire   [2:2]     RX_DATA_0_slice_28;
wire   [3:3]     RX_DATA_0_slice_29;
wire   [4:4]     RX_DATA_0_slice_30;
wire   [5:5]     RX_DATA_0_slice_31;
wire   [0:0]     RX_DATA_0_slice_32;
wire   [1:1]     RX_DATA_0_slice_33;
wire   [2:2]     RX_DATA_0_slice_34;
wire   [3:3]     RX_DATA_0_slice_35;
wire   [4:4]     RX_DATA_0_slice_36;
wire   [5:5]     RX_DATA_0_slice_37;
wire   [3:0]     TX_DATA_0_net_0;
wire   [3:0]     TX_DATA_1_net_0;
wire   [3:0]     TX_DATA_2_net_0;
wire   [3:0]     TX_DATA_3_net_0;
wire   [3:0]     TX_DATA_4_net_0;
wire   [3:0]     TX_DATA_5_net_0;
wire   [3:0]     TX_DATA_6_net_0;
wire   [3:0]     TX_DATA_7_net_0;
wire   [3:0]     TX_DATA_8_net_0;
wire   [3:0]     TX_DATA_9_net_0;
wire   [3:0]     TX_DATA_10_net_0;
wire   [3:0]     TX_DATA_11_net_0;
wire   [3:0]     TX_DATA_0_net_1;
wire   [3:0]     OE_DATA_0_net_0;
wire   [3:0]     TX_DATA_0_net_2;
wire   [3:0]     TX_DATA_0_net_3;
wire   [3:0]     TX_DATA_0_net_4;
wire   [3:0]     TX_DATA_1_net_1;
wire   [3:0]     TX_DATA_0_net_5;
wire   [3:0]     TX_DATA_1_net_2;
wire   [3:0]     TX_DATA_0_net_6;
wire   [3:0]     TX_DATA_0_net_7;
wire   [3:0]     TX_DATA_0_net_8;
wire   [3:0]     TX_DATA_0_net_9;
wire   [3:0]     TX_DATA_0_net_10;
wire   [3:0]     TX_DATA_0_net_11;
wire   [3:0]     TX_DATA_0_net_12;
wire   [1:0]     HS_IO_CLK_net_0;
wire   [2:0]     READ_CLK_SEL_net_0;
wire   [7:0]     TX_DATA_0_net_13;
wire   [3:0]     OE_DATA_0_net_1;
wire   [7:0]     TX_DATA_0_net_14;
wire   [7:0]     TX_DATA_1_net_3;
wire   [7:0]     TX_DATA_2_net_1;
wire   [7:0]     TX_DATA_3_net_1;
wire   [7:0]     TX_DATA_4_net_1;
wire   [7:0]     TX_DATA_5_net_1;
wire   [7:0]     TX_DATA_6_net_1;
wire   [7:0]     TX_DATA_7_net_1;
wire   [3:0]     OE_DATA_0_net_2;
wire   [3:0]     OE_DATA_1_net_0;
wire   [3:0]     OE_DATA_2_net_0;
wire   [3:0]     OE_DATA_3_net_0;
wire   [3:0]     OE_DATA_4_net_0;
wire   [3:0]     OE_DATA_5_net_0;
wire   [3:0]     OE_DATA_6_net_0;
wire   [3:0]     OE_DATA_7_net_0;
wire   [3:0]     OE_DATA_0_net_3;
wire   [7:0]     TX_DATA_0_net_15;
wire   [3:0]     OE_DATA_0_net_4;
wire   [1:0]     HS_IO_CLK_net_1;
wire   [2:0]     READ_CLK_SEL_net_1;
wire   [7:0]     TX_DATA_0_net_16;
wire   [3:0]     OE_DATA_0_net_5;
wire   [7:0]     TX_DATA_0_net_17;
wire   [7:0]     TX_DATA_1_net_4;
wire   [7:0]     TX_DATA_2_net_2;
wire   [7:0]     TX_DATA_3_net_2;
wire   [7:0]     TX_DATA_4_net_2;
wire   [7:0]     TX_DATA_5_net_2;
wire   [7:0]     TX_DATA_6_net_2;
wire   [7:0]     TX_DATA_7_net_2;
wire   [3:0]     OE_DATA_0_net_6;
wire   [3:0]     OE_DATA_1_net_1;
wire   [3:0]     OE_DATA_2_net_1;
wire   [3:0]     OE_DATA_3_net_1;
wire   [3:0]     OE_DATA_4_net_1;
wire   [3:0]     OE_DATA_5_net_1;
wire   [3:0]     OE_DATA_6_net_1;
wire   [3:0]     OE_DATA_7_net_1;
wire   [3:0]     OE_DATA_0_net_7;
wire   [7:0]     TX_DATA_0_net_18;
wire   [3:0]     OE_DATA_0_net_8;
wire   [1:0]     HS_IO_CLK_net_2;
wire   [2:0]     READ_CLK_SEL_net_2;
wire   [7:0]     TX_DATA_0_net_19;
wire   [3:0]     OE_DATA_0_net_9;
wire   [7:0]     TX_DATA_0_net_20;
wire   [7:0]     TX_DATA_1_net_5;
wire   [7:0]     TX_DATA_2_net_3;
wire   [7:0]     TX_DATA_3_net_3;
wire   [7:0]     TX_DATA_4_net_3;
wire   [7:0]     TX_DATA_5_net_3;
wire   [7:0]     TX_DATA_6_net_3;
wire   [7:0]     TX_DATA_7_net_3;
wire   [3:0]     OE_DATA_0_net_10;
wire   [3:0]     OE_DATA_1_net_2;
wire   [3:0]     OE_DATA_2_net_2;
wire   [3:0]     OE_DATA_3_net_2;
wire   [3:0]     OE_DATA_4_net_2;
wire   [3:0]     OE_DATA_5_net_2;
wire   [3:0]     OE_DATA_6_net_2;
wire   [3:0]     OE_DATA_7_net_2;
wire   [3:0]     OE_DATA_0_net_11;
wire   [7:0]     TX_DATA_0_net_21;
wire   [3:0]     OE_DATA_0_net_12;
wire   [1:0]     HS_IO_CLK_net_3;
wire   [2:0]     READ_CLK_SEL_net_3;
wire   [7:0]     TX_DATA_0_net_22;
wire   [3:0]     OE_DATA_0_net_13;
wire   [7:0]     TX_DATA_0_net_23;
wire   [7:0]     TX_DATA_1_net_6;
wire   [7:0]     TX_DATA_2_net_4;
wire   [7:0]     TX_DATA_3_net_4;
wire   [7:0]     TX_DATA_4_net_4;
wire   [7:0]     TX_DATA_5_net_4;
wire   [7:0]     TX_DATA_6_net_4;
wire   [7:0]     TX_DATA_7_net_4;
wire   [3:0]     OE_DATA_0_net_14;
wire   [3:0]     OE_DATA_1_net_3;
wire   [3:0]     OE_DATA_2_net_3;
wire   [3:0]     OE_DATA_3_net_3;
wire   [3:0]     OE_DATA_4_net_3;
wire   [3:0]     OE_DATA_5_net_3;
wire   [3:0]     OE_DATA_6_net_3;
wire   [3:0]     OE_DATA_7_net_3;
wire   [3:0]     OE_DATA_0_net_15;
wire   [7:0]     TX_DATA_0_net_24;
wire   [3:0]     OE_DATA_0_net_16;
wire   [16:0]    DFI_ADDRESS_P0;
wire   [1:0]     DFI_BG_P0;
wire   [1:0]     DFI_BANK_P0;
wire   [16:0]    DFI_ADDRESS_P1;
wire   [1:0]     DFI_BG_P1;
wire   [1:0]     DFI_BANK_P1;
wire   [16:0]    DFI_ADDRESS_P2;
wire   [1:0]     DFI_BG_P2;
wire   [1:0]     DFI_BANK_P2;
wire   [16:0]    DFI_ADDRESS_P3;
wire   [1:0]     DFI_BG_P3;
wire   [1:0]     DFI_BANK_P3;
wire   [31:0]    DFI_WRDATA_EN_P0;
wire   [7:0]     DFI_WRDATA_MASK_P0;
wire   [63:0]    DFI_WRDATA_P0;
wire   [31:0]    DFI_WRDATA_EN_P1;
wire   [7:0]     DFI_WRDATA_MASK_P1;
wire   [63:0]    DFI_WRDATA_P1;
wire   [31:0]    DFI_WRDATA_EN_P2;
wire   [7:0]     DFI_WRDATA_MASK_P2;
wire   [63:0]    DFI_WRDATA_P2;
wire   [31:0]    DFI_WRDATA_EN_P3;
wire   [7:0]     DFI_WRDATA_MASK_P3;
wire   [63:0]    DFI_WRDATA_P3;
wire   [31:0]    DFI_RDDATA_EN_P0;
wire   [31:0]    DFI_RDDATA_EN_P1;
wire   [31:0]    DFI_RDDATA_EN_P2;
wire   [31:0]    DFI_RDDATA_EN_P3;
wire   [11:0]    PAD_O_net_0;
wire   [3:0]     RX_DATA_0_net_0;
wire   [7:0]     RX_DATA_0_net_1;
wire   [7:0]     RX_DATA_0_net_2;
wire   [3:0]     BURST_DETECT_net_0;
wire   [11:0]    CLK_SEL_net_0;
wire   [3:0]     DELAY_LINE_SEL_RD_net_0;
wire   [35:0]    DIRECTION_net_0;
wire   [3:0]     IOG_OE_P0_net_0;
wire   [3:0]     IOG_OE_P1_net_0;
wire   [3:0]     IOG_OE_P2_net_0;
wire   [3:0]     IOG_OE_P3_net_0;
wire   [3:0]     DQS_OE_P0_net_0;
wire   [3:0]     DQS_OE_P1_net_0;
wire   [3:0]     DQS_OE_P2_net_0;
wire   [3:0]     DQS_OE_P3_net_0;
wire   [3:0]     DM_OE_P0_net_0;
wire   [3:0]     DM_OE_P1_net_0;
wire   [3:0]     DM_OE_P2_net_0;
wire   [3:0]     DM_OE_P3_net_0;
wire   [35:0]    LOAD_net_0;
wire   [35:0]    MOVE_net_0;
wire   [35:0]    RX_OUT_OF_RANGE_net_0;
wire   [35:0]    TX_OUT_OF_RANGE_net_0;
wire   [3:0]     ODT_DYN_LANE_net_0;
wire   [255:0]   IOG_RDDATA_net_0;
wire   [3:0]     IOG_RDDATA_VALID_net_0;
wire   [31:0]    PAD_RDDATA_net_0;
wire   [3:0]     IOG_RDDATA_EN_P0_P_net_0;
wire   [3:0]     IOG_RDDATA_EN_P0_N_net_0;
wire   [3:0]     IOG_RDDATA_EN_P1_P_net_0;
wire   [3:0]     IOG_RDDATA_EN_P1_N_net_0;
wire   [3:0]     IOG_RDDATA_EN_P2_P_net_0;
wire   [3:0]     IOG_RDDATA_EN_P2_N_net_0;
wire   [3:0]     IOG_RDDATA_EN_P3_P_net_0;
wire   [3:0]     IOG_RDDATA_EN_P3_N_net_0;
wire   [3:0]     DQSW_EYE_MONITOR_CLR_FLAGS_net_0;
wire   [3:0]     DQSW_EYE_MONITOR_EARLY_net_0;
wire   [3:0]     DQSW_EYE_MONITOR_LATE_net_0;
wire   [3:0]     DQSW270_EYE_MONITOR_CLR_FLAGS_net_0;
wire   [3:0]     DQSW270_EYE_MONITOR_EARLY_net_0;
wire   [3:0]     DQSW270_EYE_MONITOR_LATE_net_0;
wire   [3:0]     DQSW_DELAY_LINE_LOAD_net_0;
wire   [3:0]     DQSW_DELAY_LINE_MOVE_net_0;
wire   [3:0]     DQSW_DELAY_LINE_DIRECTION_net_0;
wire   [3:0]     DQSW270_DELAY_LINE_LOAD_net_0;
wire   [3:0]     DQSW270_DELAY_LINE_MOVE_net_0;
wire   [3:0]     DQSW270_DELAY_LINE_DIRECTION_net_0;
wire   [31:0]    DQSW_SELA_net_0;
wire   [3:0]     DQSW270_IGEAR_RX8_net_0;
wire   [3:0]     DQSW_DELAY_LINE_OOR_net_0;
wire   [3:0]     DQSW270_DELAY_LINE_OOR_net_0;
wire   [3:0]     INIT_PAUSE_net_0;
wire   [19:0]    DFI_ADDRESS_P0_net_0;
wire   [19:0]    DFI_ADDRESS_P1_net_0;
wire   [19:0]    DFI_ADDRESS_P2_net_0;
wire   [19:0]    DFI_ADDRESS_P3_net_0;
wire   [7:0]     IOG_WRDATA_MASK_P0_net_0;
wire   [7:0]     IOG_WRDATA_MASK_P1_net_0;
wire   [7:0]     IOG_WRDATA_MASK_P2_net_0;
wire   [7:0]     IOG_WRDATA_MASK_P3_net_0;
wire   [19:0]    IOG_ADDRESS_P0_net_0;
wire   [19:0]    IOG_ADDRESS_P1_net_0;
wire   [19:0]    IOG_ADDRESS_P2_net_0;
wire   [19:0]    IOG_ADDRESS_P3_net_0;
wire   [3:0]     BCLK_IGEAR_RX_net_0;
wire   [7:0]     DQSW270_IGEAR_RX_net_0;
wire   [7:0]     DQSW_IGEAR_RX_net_0;
wire   [255:0]   IOG_DQ_TXDATA_IN_net_0;
wire   [255:0]   IOG_DQ_TXDATA_OUT_net_0;
wire   [31:0]    IOG_DM_TXDATA_IN_net_0;
wire   [31:0]    IOG_DM_TXDATA_OUT_net_0;
wire   [3:0]     DFI_BANK_P0_net_0;
wire   [3:0]     DFI_BANK_P1_net_0;
wire   [3:0]     DFI_BANK_P2_net_0;
wire   [3:0]     DFI_BANK_P3_net_0;
wire   [3:0]     DFI_BANK_P0_OUT_net_0;
wire   [3:0]     DFI_BANK_P1_OUT_net_0;
wire   [3:0]     DFI_BANK_P2_OUT_net_0;
wire   [3:0]     DFI_BANK_P3_OUT_net_0;
wire   [1:0]     DFI_BG_P0_net_0;
wire   [1:0]     DFI_BG_P1_net_0;
wire   [1:0]     DFI_BG_P2_net_0;
wire   [1:0]     DFI_BG_P3_net_0;
wire   [1:0]     DFI_BG_P0_OUT_net_0;
wire   [1:0]     DFI_BG_P1_OUT_net_0;
wire   [1:0]     DFI_BG_P2_OUT_net_0;
wire   [1:0]     DFI_BG_P3_OUT_net_0;
wire   [7:0]     RX_DATA_0_net_3;
wire   [7:0]     RX_DATA_1_net_0;
wire   [7:0]     RX_DATA_2_net_0;
wire   [7:0]     RX_DATA_3_net_0;
wire   [7:0]     RX_DATA_4_net_0;
wire   [7:0]     RX_DATA_5_net_0;
wire   [7:0]     RX_DATA_6_net_0;
wire   [7:0]     RX_DATA_7_net_0;
wire   [7:0]     PAD_net_0;
wire   [1:0]     RX_DATA_0_net_4;
wire   [7:0]     RX_DATA_0_net_5;
wire   [7:0]     RX_DATA_0_net_6;
wire   [7:0]     RX_DATA_1_net_1;
wire   [7:0]     RX_DATA_2_net_1;
wire   [7:0]     RX_DATA_3_net_1;
wire   [7:0]     RX_DATA_4_net_1;
wire   [7:0]     RX_DATA_5_net_1;
wire   [7:0]     RX_DATA_6_net_1;
wire   [7:0]     RX_DATA_7_net_1;
wire   [7:0]     PAD_net_1;
wire   [1:0]     RX_DATA_0_net_7;
wire   [7:0]     RX_DATA_0_net_8;
wire   [7:0]     RX_DATA_0_net_9;
wire   [7:0]     RX_DATA_1_net_2;
wire   [7:0]     RX_DATA_2_net_2;
wire   [7:0]     RX_DATA_3_net_2;
wire   [7:0]     RX_DATA_4_net_2;
wire   [7:0]     RX_DATA_5_net_2;
wire   [7:0]     RX_DATA_6_net_2;
wire   [7:0]     RX_DATA_7_net_2;
wire   [7:0]     PAD_net_2;
wire   [1:0]     RX_DATA_0_net_10;
wire   [7:0]     RX_DATA_0_net_11;
wire   [7:0]     RX_DATA_0_net_12;
wire   [7:0]     RX_DATA_1_net_3;
wire   [7:0]     RX_DATA_2_net_3;
wire   [7:0]     RX_DATA_3_net_3;
wire   [7:0]     RX_DATA_4_net_3;
wire   [7:0]     RX_DATA_5_net_3;
wire   [7:0]     RX_DATA_6_net_3;
wire   [7:0]     RX_DATA_7_net_3;
wire   [7:0]     PAD_net_3;
wire   [1:0]     RX_DATA_0_net_13;
wire   [7:0]     RX_DATA_0_net_14;
//--------------------------------------------------------------------
// TiedOff Nets
//--------------------------------------------------------------------
wire   [1:0]     DFI_CALVL_RESP_const_net_0;
wire             VCC_net;
wire             GND_net;
wire   [1:0]     DFI_PHYUPD_TYPE_const_net_0;
wire   [3:0]     OE_DATA_0_const_net_0;
wire   [3:0]     OE_DATA_1_const_net_0;
wire   [3:0]     OE_DATA_2_const_net_0;
wire   [3:0]     OE_DATA_3_const_net_0;
wire   [3:0]     OE_DATA_4_const_net_0;
wire   [3:0]     OE_DATA_5_const_net_0;
wire   [3:0]     OE_DATA_6_const_net_0;
wire   [3:0]     OE_DATA_7_const_net_0;
wire   [3:0]     OE_DATA_8_const_net_0;
wire   [3:0]     OE_DATA_9_const_net_0;
wire   [3:0]     OE_DATA_10_const_net_0;
wire   [3:0]     OE_DATA_11_const_net_0;
wire   [3:0]     OE_DATA_0_const_net_1;
wire   [3:0]     OE_DATA_0_const_net_2;
wire   [3:0]     OE_DATA_0_const_net_3;
wire   [3:0]     OE_DATA_1_const_net_1;
wire   [3:0]     OE_DATA_0_const_net_4;
wire   [3:0]     OE_DATA_1_const_net_2;
wire   [3:0]     OE_DATA_0_const_net_5;
wire   [3:0]     OE_DATA_0_const_net_6;
wire   [3:0]     OE_DATA_0_const_net_7;
wire   [3:0]     OE_DATA_0_const_net_8;
wire   [3:0]     OE_DATA_0_const_net_9;
wire   [3:0]     OE_DATA_0_const_net_10;
wire   [7:0]     TRAINING_PATTERN_const_net_0;
wire   [3:0]     OE_DATA_0_const_net_11;
wire   [2:0]     EYE_MONITOR_WIDTH_IN_const_net_0;
wire   [7:0]     TX_DATA_0_const_net_0;
wire   [1:0]     TX_DATA_0_const_net_1;
wire   [1:0]     OE_DATA_0_const_net_12;
wire   [2:0]     EYE_MONITOR_WIDTH_IN_const_net_1;
wire   [7:0]     TX_DATA_0_const_net_2;
wire   [1:0]     TX_DATA_0_const_net_3;
wire   [1:0]     OE_DATA_0_const_net_13;
wire   [2:0]     EYE_MONITOR_WIDTH_IN_const_net_2;
wire   [7:0]     TX_DATA_0_const_net_4;
wire   [1:0]     TX_DATA_0_const_net_5;
wire   [1:0]     OE_DATA_0_const_net_14;
wire   [2:0]     EYE_MONITOR_WIDTH_IN_const_net_3;
wire   [7:0]     TX_DATA_0_const_net_6;
wire   [1:0]     TX_DATA_0_const_net_7;
wire   [1:0]     OE_DATA_0_const_net_15;
wire   [1:0]     RX_DQS_90_const_net_0;
wire   [2:0]     FIFO_WR_PTR_const_net_0;
wire   [2:0]     FIFO_RD_PTR_const_net_0;
wire   [2:0]     EYE_MONITOR_LANE_WIDTH_const_net_0;
wire   [3:0]     TX_DATA_12_const_net_0;
wire   [3:0]     TX_DATA_13_const_net_0;
wire   [3:0]     TX_DATA_14_const_net_0;
wire   [3:0]     TX_DATA_15_const_net_0;
wire   [3:0]     TX_DATA_16_const_net_0;
wire   [3:0]     TX_DATA_17_const_net_0;
wire   [3:0]     TX_DATA_18_const_net_0;
wire   [3:0]     TX_DATA_19_const_net_0;
wire   [3:0]     TX_DATA_20_const_net_0;
wire   [3:0]     TX_DATA_21_const_net_0;
wire   [3:0]     TX_DATA_22_const_net_0;
wire   [3:0]     TX_DATA_23_const_net_0;
wire   [3:0]     TX_DATA_24_const_net_0;
wire   [3:0]     TX_DATA_25_const_net_0;
wire   [3:0]     TX_DATA_26_const_net_0;
wire   [3:0]     TX_DATA_27_const_net_0;
wire   [3:0]     TX_DATA_28_const_net_0;
wire   [3:0]     TX_DATA_29_const_net_0;
wire   [3:0]     TX_DATA_30_const_net_0;
wire   [3:0]     TX_DATA_31_const_net_0;
wire   [3:0]     TX_DATA_32_const_net_0;
wire   [3:0]     TX_DATA_33_const_net_0;
wire   [3:0]     TX_DATA_34_const_net_0;
wire   [3:0]     TX_DATA_35_const_net_0;
wire   [3:0]     TX_DATA_36_const_net_0;
wire   [3:0]     TX_DATA_37_const_net_0;
wire   [3:0]     TX_DATA_38_const_net_0;
wire   [3:0]     TX_DATA_39_const_net_0;
wire   [3:0]     TX_DATA_40_const_net_0;
wire   [3:0]     TX_DATA_41_const_net_0;
wire   [3:0]     TX_DATA_42_const_net_0;
wire   [3:0]     TX_DATA_43_const_net_0;
wire   [3:0]     TX_DATA_44_const_net_0;
wire   [3:0]     TX_DATA_45_const_net_0;
wire   [3:0]     TX_DATA_46_const_net_0;
wire   [3:0]     TX_DATA_47_const_net_0;
wire   [3:0]     TX_DATA_48_const_net_0;
wire   [3:0]     TX_DATA_49_const_net_0;
wire   [3:0]     TX_DATA_50_const_net_0;
wire   [3:0]     TX_DATA_51_const_net_0;
wire   [3:0]     TX_DATA_52_const_net_0;
wire   [3:0]     TX_DATA_53_const_net_0;
wire   [3:0]     TX_DATA_54_const_net_0;
wire   [3:0]     TX_DATA_55_const_net_0;
wire   [3:0]     TX_DATA_56_const_net_0;
wire   [3:0]     TX_DATA_57_const_net_0;
wire   [3:0]     TX_DATA_58_const_net_0;
wire   [3:0]     TX_DATA_59_const_net_0;
wire   [3:0]     TX_DATA_60_const_net_0;
wire   [3:0]     TX_DATA_61_const_net_0;
wire   [3:0]     TX_DATA_62_const_net_0;
wire   [3:0]     TX_DATA_63_const_net_0;
wire   [3:0]     TX_DATA_64_const_net_0;
wire   [3:0]     TX_DATA_65_const_net_0;
wire   [3:0]     TX_DATA_66_const_net_0;
wire   [3:0]     TX_DATA_67_const_net_0;
wire   [3:0]     TX_DATA_68_const_net_0;
wire   [3:0]     TX_DATA_69_const_net_0;
wire   [3:0]     TX_DATA_70_const_net_0;
wire   [3:0]     TX_DATA_71_const_net_0;
wire   [3:0]     TX_DATA_72_const_net_0;
wire   [3:0]     TX_DATA_73_const_net_0;
wire   [3:0]     TX_DATA_74_const_net_0;
wire   [3:0]     TX_DATA_75_const_net_0;
wire   [3:0]     TX_DATA_76_const_net_0;
wire   [3:0]     TX_DATA_77_const_net_0;
wire   [3:0]     TX_DATA_78_const_net_0;
wire   [3:0]     TX_DATA_79_const_net_0;
wire   [3:0]     TX_DATA_80_const_net_0;
wire   [3:0]     TX_DATA_81_const_net_0;
wire   [3:0]     TX_DATA_82_const_net_0;
wire   [3:0]     TX_DATA_83_const_net_0;
wire   [3:0]     TX_DATA_84_const_net_0;
wire   [3:0]     TX_DATA_85_const_net_0;
wire   [3:0]     TX_DATA_86_const_net_0;
wire   [3:0]     TX_DATA_87_const_net_0;
wire   [3:0]     TX_DATA_88_const_net_0;
wire   [3:0]     TX_DATA_89_const_net_0;
wire   [3:0]     TX_DATA_90_const_net_0;
wire   [3:0]     TX_DATA_91_const_net_0;
wire   [3:0]     TX_DATA_92_const_net_0;
wire   [3:0]     TX_DATA_93_const_net_0;
wire   [3:0]     TX_DATA_94_const_net_0;
wire   [3:0]     TX_DATA_95_const_net_0;
wire   [3:0]     TX_DATA_96_const_net_0;
wire   [3:0]     TX_DATA_97_const_net_0;
wire   [3:0]     TX_DATA_98_const_net_0;
wire   [3:0]     TX_DATA_99_const_net_0;
wire   [3:0]     TX_DATA_100_const_net_0;
wire   [3:0]     TX_DATA_101_const_net_0;
wire   [3:0]     TX_DATA_102_const_net_0;
wire   [3:0]     TX_DATA_103_const_net_0;
wire   [3:0]     TX_DATA_104_const_net_0;
wire   [3:0]     TX_DATA_105_const_net_0;
wire   [3:0]     TX_DATA_106_const_net_0;
wire   [3:0]     TX_DATA_107_const_net_0;
wire   [3:0]     TX_DATA_108_const_net_0;
wire   [3:0]     TX_DATA_109_const_net_0;
wire   [3:0]     TX_DATA_110_const_net_0;
wire   [3:0]     TX_DATA_111_const_net_0;
wire   [3:0]     TX_DATA_112_const_net_0;
wire   [3:0]     TX_DATA_113_const_net_0;
wire   [3:0]     TX_DATA_114_const_net_0;
wire   [3:0]     TX_DATA_115_const_net_0;
wire   [3:0]     TX_DATA_116_const_net_0;
wire   [3:0]     TX_DATA_117_const_net_0;
wire   [3:0]     TX_DATA_118_const_net_0;
wire   [3:0]     TX_DATA_119_const_net_0;
wire   [3:0]     TX_DATA_120_const_net_0;
wire   [3:0]     TX_DATA_121_const_net_0;
wire   [3:0]     TX_DATA_122_const_net_0;
wire   [3:0]     TX_DATA_123_const_net_0;
wire   [3:0]     TX_DATA_124_const_net_0;
wire   [3:0]     TX_DATA_125_const_net_0;
wire   [3:0]     TX_DATA_126_const_net_0;
wire   [3:0]     TX_DATA_127_const_net_0;
wire   [3:0]     OE_DATA_12_const_net_0;
wire   [3:0]     OE_DATA_13_const_net_0;
wire   [3:0]     OE_DATA_14_const_net_0;
wire   [3:0]     OE_DATA_15_const_net_0;
wire   [3:0]     OE_DATA_16_const_net_0;
wire   [3:0]     OE_DATA_17_const_net_0;
wire   [3:0]     OE_DATA_18_const_net_0;
wire   [3:0]     OE_DATA_19_const_net_0;
wire   [3:0]     OE_DATA_20_const_net_0;
wire   [3:0]     OE_DATA_21_const_net_0;
wire   [3:0]     OE_DATA_22_const_net_0;
wire   [3:0]     OE_DATA_23_const_net_0;
wire   [3:0]     OE_DATA_24_const_net_0;
wire   [3:0]     OE_DATA_25_const_net_0;
wire   [3:0]     OE_DATA_26_const_net_0;
wire   [3:0]     OE_DATA_27_const_net_0;
wire   [3:0]     OE_DATA_28_const_net_0;
wire   [3:0]     OE_DATA_29_const_net_0;
wire   [3:0]     OE_DATA_30_const_net_0;
wire   [3:0]     OE_DATA_31_const_net_0;
wire   [3:0]     OE_DATA_32_const_net_0;
wire   [3:0]     OE_DATA_33_const_net_0;
wire   [3:0]     OE_DATA_34_const_net_0;
wire   [3:0]     OE_DATA_35_const_net_0;
wire   [3:0]     OE_DATA_36_const_net_0;
wire   [3:0]     OE_DATA_37_const_net_0;
wire   [3:0]     OE_DATA_38_const_net_0;
wire   [3:0]     OE_DATA_39_const_net_0;
wire   [3:0]     OE_DATA_40_const_net_0;
wire   [3:0]     OE_DATA_41_const_net_0;
wire   [3:0]     OE_DATA_42_const_net_0;
wire   [3:0]     OE_DATA_43_const_net_0;
wire   [3:0]     OE_DATA_44_const_net_0;
wire   [3:0]     OE_DATA_45_const_net_0;
wire   [3:0]     OE_DATA_46_const_net_0;
wire   [3:0]     OE_DATA_47_const_net_0;
wire   [3:0]     OE_DATA_48_const_net_0;
wire   [3:0]     OE_DATA_49_const_net_0;
wire   [3:0]     OE_DATA_50_const_net_0;
wire   [3:0]     OE_DATA_51_const_net_0;
wire   [3:0]     OE_DATA_52_const_net_0;
wire   [3:0]     OE_DATA_53_const_net_0;
wire   [3:0]     OE_DATA_54_const_net_0;
wire   [3:0]     OE_DATA_55_const_net_0;
wire   [3:0]     OE_DATA_56_const_net_0;
wire   [3:0]     OE_DATA_57_const_net_0;
wire   [3:0]     OE_DATA_58_const_net_0;
wire   [3:0]     OE_DATA_59_const_net_0;
wire   [3:0]     OE_DATA_60_const_net_0;
wire   [3:0]     OE_DATA_61_const_net_0;
wire   [3:0]     OE_DATA_62_const_net_0;
wire   [3:0]     OE_DATA_63_const_net_0;
wire   [3:0]     OE_DATA_64_const_net_0;
wire   [3:0]     OE_DATA_65_const_net_0;
wire   [3:0]     OE_DATA_66_const_net_0;
wire   [3:0]     OE_DATA_67_const_net_0;
wire   [3:0]     OE_DATA_68_const_net_0;
wire   [3:0]     OE_DATA_69_const_net_0;
wire   [3:0]     OE_DATA_70_const_net_0;
wire   [3:0]     OE_DATA_71_const_net_0;
wire   [3:0]     OE_DATA_72_const_net_0;
wire   [3:0]     OE_DATA_73_const_net_0;
wire   [3:0]     OE_DATA_74_const_net_0;
wire   [3:0]     OE_DATA_75_const_net_0;
wire   [3:0]     OE_DATA_76_const_net_0;
wire   [3:0]     OE_DATA_77_const_net_0;
wire   [3:0]     OE_DATA_78_const_net_0;
wire   [3:0]     OE_DATA_79_const_net_0;
wire   [3:0]     OE_DATA_80_const_net_0;
wire   [3:0]     OE_DATA_81_const_net_0;
wire   [3:0]     OE_DATA_82_const_net_0;
wire   [3:0]     OE_DATA_83_const_net_0;
wire   [3:0]     OE_DATA_84_const_net_0;
wire   [3:0]     OE_DATA_85_const_net_0;
wire   [3:0]     OE_DATA_86_const_net_0;
wire   [3:0]     OE_DATA_87_const_net_0;
wire   [3:0]     OE_DATA_88_const_net_0;
wire   [3:0]     OE_DATA_89_const_net_0;
wire   [3:0]     OE_DATA_90_const_net_0;
wire   [3:0]     OE_DATA_91_const_net_0;
wire   [3:0]     OE_DATA_92_const_net_0;
wire   [3:0]     OE_DATA_93_const_net_0;
wire   [3:0]     OE_DATA_94_const_net_0;
wire   [3:0]     OE_DATA_95_const_net_0;
wire   [3:0]     OE_DATA_96_const_net_0;
wire   [3:0]     OE_DATA_97_const_net_0;
wire   [3:0]     OE_DATA_98_const_net_0;
wire   [3:0]     OE_DATA_99_const_net_0;
wire   [3:0]     OE_DATA_100_const_net_0;
wire   [3:0]     OE_DATA_101_const_net_0;
wire   [3:0]     OE_DATA_102_const_net_0;
wire   [3:0]     OE_DATA_103_const_net_0;
wire   [3:0]     OE_DATA_104_const_net_0;
wire   [3:0]     OE_DATA_105_const_net_0;
wire   [3:0]     OE_DATA_106_const_net_0;
wire   [3:0]     OE_DATA_107_const_net_0;
wire   [3:0]     OE_DATA_108_const_net_0;
wire   [3:0]     OE_DATA_109_const_net_0;
wire   [3:0]     OE_DATA_110_const_net_0;
wire   [3:0]     OE_DATA_111_const_net_0;
wire   [3:0]     OE_DATA_112_const_net_0;
wire   [3:0]     OE_DATA_113_const_net_0;
wire   [3:0]     OE_DATA_114_const_net_0;
wire   [3:0]     OE_DATA_115_const_net_0;
wire   [3:0]     OE_DATA_116_const_net_0;
wire   [3:0]     OE_DATA_117_const_net_0;
wire   [3:0]     OE_DATA_118_const_net_0;
wire   [3:0]     OE_DATA_119_const_net_0;
wire   [3:0]     OE_DATA_120_const_net_0;
wire   [3:0]     OE_DATA_121_const_net_0;
wire   [3:0]     OE_DATA_122_const_net_0;
wire   [3:0]     OE_DATA_123_const_net_0;
wire   [3:0]     OE_DATA_124_const_net_0;
wire   [3:0]     OE_DATA_125_const_net_0;
wire   [3:0]     OE_DATA_126_const_net_0;
wire   [3:0]     OE_DATA_127_const_net_0;
wire   [11:0]    PAD_const_net_0;
wire   [11:0]    PAD_I_const_net_0;
wire   [11:0]    PAD_N_const_net_0;
wire   [11:0]    PAD_I_N_const_net_0;
wire   [1:0]     RX_DQS_90_const_net_1;
wire   [2:0]     FIFO_WR_PTR_const_net_1;
wire   [2:0]     FIFO_RD_PTR_const_net_1;
wire   [2:0]     EYE_MONITOR_LANE_WIDTH_const_net_1;
wire   [3:0]     TX_DATA_1_const_net_0;
wire   [3:0]     TX_DATA_2_const_net_0;
wire   [3:0]     TX_DATA_3_const_net_0;
wire   [3:0]     TX_DATA_4_const_net_0;
wire   [3:0]     TX_DATA_5_const_net_0;
wire   [3:0]     TX_DATA_6_const_net_0;
wire   [3:0]     TX_DATA_7_const_net_0;
wire   [3:0]     TX_DATA_8_const_net_0;
wire   [3:0]     TX_DATA_9_const_net_0;
wire   [3:0]     TX_DATA_10_const_net_0;
wire   [3:0]     TX_DATA_11_const_net_0;
wire   [3:0]     TX_DATA_12_const_net_1;
wire   [3:0]     TX_DATA_13_const_net_1;
wire   [3:0]     TX_DATA_14_const_net_1;
wire   [3:0]     TX_DATA_15_const_net_1;
wire   [3:0]     TX_DATA_16_const_net_1;
wire   [3:0]     TX_DATA_17_const_net_1;
wire   [3:0]     TX_DATA_18_const_net_1;
wire   [3:0]     TX_DATA_19_const_net_1;
wire   [3:0]     TX_DATA_20_const_net_1;
wire   [3:0]     TX_DATA_21_const_net_1;
wire   [3:0]     TX_DATA_22_const_net_1;
wire   [3:0]     TX_DATA_23_const_net_1;
wire   [3:0]     TX_DATA_24_const_net_1;
wire   [3:0]     TX_DATA_25_const_net_1;
wire   [3:0]     TX_DATA_26_const_net_1;
wire   [3:0]     TX_DATA_27_const_net_1;
wire   [3:0]     TX_DATA_28_const_net_1;
wire   [3:0]     TX_DATA_29_const_net_1;
wire   [3:0]     TX_DATA_30_const_net_1;
wire   [3:0]     TX_DATA_31_const_net_1;
wire   [3:0]     TX_DATA_32_const_net_1;
wire   [3:0]     TX_DATA_33_const_net_1;
wire   [3:0]     TX_DATA_34_const_net_1;
wire   [3:0]     TX_DATA_35_const_net_1;
wire   [3:0]     TX_DATA_36_const_net_1;
wire   [3:0]     TX_DATA_37_const_net_1;
wire   [3:0]     TX_DATA_38_const_net_1;
wire   [3:0]     TX_DATA_39_const_net_1;
wire   [3:0]     TX_DATA_40_const_net_1;
wire   [3:0]     TX_DATA_41_const_net_1;
wire   [3:0]     TX_DATA_42_const_net_1;
wire   [3:0]     TX_DATA_43_const_net_1;
wire   [3:0]     TX_DATA_44_const_net_1;
wire   [3:0]     TX_DATA_45_const_net_1;
wire   [3:0]     TX_DATA_46_const_net_1;
wire   [3:0]     TX_DATA_47_const_net_1;
wire   [3:0]     TX_DATA_48_const_net_1;
wire   [3:0]     TX_DATA_49_const_net_1;
wire   [3:0]     TX_DATA_50_const_net_1;
wire   [3:0]     TX_DATA_51_const_net_1;
wire   [3:0]     TX_DATA_52_const_net_1;
wire   [3:0]     TX_DATA_53_const_net_1;
wire   [3:0]     TX_DATA_54_const_net_1;
wire   [3:0]     TX_DATA_55_const_net_1;
wire   [3:0]     TX_DATA_56_const_net_1;
wire   [3:0]     TX_DATA_57_const_net_1;
wire   [3:0]     TX_DATA_58_const_net_1;
wire   [3:0]     TX_DATA_59_const_net_1;
wire   [3:0]     TX_DATA_60_const_net_1;
wire   [3:0]     TX_DATA_61_const_net_1;
wire   [3:0]     TX_DATA_62_const_net_1;
wire   [3:0]     TX_DATA_63_const_net_1;
wire   [3:0]     TX_DATA_64_const_net_1;
wire   [3:0]     TX_DATA_65_const_net_1;
wire   [3:0]     TX_DATA_66_const_net_1;
wire   [3:0]     TX_DATA_67_const_net_1;
wire   [3:0]     TX_DATA_68_const_net_1;
wire   [3:0]     TX_DATA_69_const_net_1;
wire   [3:0]     TX_DATA_70_const_net_1;
wire   [3:0]     TX_DATA_71_const_net_1;
wire   [3:0]     TX_DATA_72_const_net_1;
wire   [3:0]     TX_DATA_73_const_net_1;
wire   [3:0]     TX_DATA_74_const_net_1;
wire   [3:0]     TX_DATA_75_const_net_1;
wire   [3:0]     TX_DATA_76_const_net_1;
wire   [3:0]     TX_DATA_77_const_net_1;
wire   [3:0]     TX_DATA_78_const_net_1;
wire   [3:0]     TX_DATA_79_const_net_1;
wire   [3:0]     TX_DATA_80_const_net_1;
wire   [3:0]     TX_DATA_81_const_net_1;
wire   [3:0]     TX_DATA_82_const_net_1;
wire   [3:0]     TX_DATA_83_const_net_1;
wire   [3:0]     TX_DATA_84_const_net_1;
wire   [3:0]     TX_DATA_85_const_net_1;
wire   [3:0]     TX_DATA_86_const_net_1;
wire   [3:0]     TX_DATA_87_const_net_1;
wire   [3:0]     TX_DATA_88_const_net_1;
wire   [3:0]     TX_DATA_89_const_net_1;
wire   [3:0]     TX_DATA_90_const_net_1;
wire   [3:0]     TX_DATA_91_const_net_1;
wire   [3:0]     TX_DATA_92_const_net_1;
wire   [3:0]     TX_DATA_93_const_net_1;
wire   [3:0]     TX_DATA_94_const_net_1;
wire   [3:0]     TX_DATA_95_const_net_1;
wire   [3:0]     TX_DATA_96_const_net_1;
wire   [3:0]     TX_DATA_97_const_net_1;
wire   [3:0]     TX_DATA_98_const_net_1;
wire   [3:0]     TX_DATA_99_const_net_1;
wire   [3:0]     TX_DATA_100_const_net_1;
wire   [3:0]     TX_DATA_101_const_net_1;
wire   [3:0]     TX_DATA_102_const_net_1;
wire   [3:0]     TX_DATA_103_const_net_1;
wire   [3:0]     TX_DATA_104_const_net_1;
wire   [3:0]     TX_DATA_105_const_net_1;
wire   [3:0]     TX_DATA_106_const_net_1;
wire   [3:0]     TX_DATA_107_const_net_1;
wire   [3:0]     TX_DATA_108_const_net_1;
wire   [3:0]     TX_DATA_109_const_net_1;
wire   [3:0]     TX_DATA_110_const_net_1;
wire   [3:0]     TX_DATA_111_const_net_1;
wire   [3:0]     TX_DATA_112_const_net_1;
wire   [3:0]     TX_DATA_113_const_net_1;
wire   [3:0]     TX_DATA_114_const_net_1;
wire   [3:0]     TX_DATA_115_const_net_1;
wire   [3:0]     TX_DATA_116_const_net_1;
wire   [3:0]     TX_DATA_117_const_net_1;
wire   [3:0]     TX_DATA_118_const_net_1;
wire   [3:0]     TX_DATA_119_const_net_1;
wire   [3:0]     TX_DATA_120_const_net_1;
wire   [3:0]     TX_DATA_121_const_net_1;
wire   [3:0]     TX_DATA_122_const_net_1;
wire   [3:0]     TX_DATA_123_const_net_1;
wire   [3:0]     TX_DATA_124_const_net_1;
wire   [3:0]     TX_DATA_125_const_net_1;
wire   [3:0]     TX_DATA_126_const_net_1;
wire   [3:0]     TX_DATA_127_const_net_1;
wire   [3:0]     OE_DATA_1_const_net_3;
wire   [3:0]     OE_DATA_2_const_net_1;
wire   [3:0]     OE_DATA_3_const_net_1;
wire   [3:0]     OE_DATA_4_const_net_1;
wire   [3:0]     OE_DATA_5_const_net_1;
wire   [3:0]     OE_DATA_6_const_net_1;
wire   [3:0]     OE_DATA_7_const_net_1;
wire   [3:0]     OE_DATA_8_const_net_1;
wire   [3:0]     OE_DATA_9_const_net_1;
wire   [3:0]     OE_DATA_10_const_net_1;
wire   [3:0]     OE_DATA_11_const_net_1;
wire   [3:0]     OE_DATA_12_const_net_1;
wire   [3:0]     OE_DATA_13_const_net_1;
wire   [3:0]     OE_DATA_14_const_net_1;
wire   [3:0]     OE_DATA_15_const_net_1;
wire   [3:0]     OE_DATA_16_const_net_1;
wire   [3:0]     OE_DATA_17_const_net_1;
wire   [3:0]     OE_DATA_18_const_net_1;
wire   [3:0]     OE_DATA_19_const_net_1;
wire   [3:0]     OE_DATA_20_const_net_1;
wire   [3:0]     OE_DATA_21_const_net_1;
wire   [3:0]     OE_DATA_22_const_net_1;
wire   [3:0]     OE_DATA_23_const_net_1;
wire   [3:0]     OE_DATA_24_const_net_1;
wire   [3:0]     OE_DATA_25_const_net_1;
wire   [3:0]     OE_DATA_26_const_net_1;
wire   [3:0]     OE_DATA_27_const_net_1;
wire   [3:0]     OE_DATA_28_const_net_1;
wire   [3:0]     OE_DATA_29_const_net_1;
wire   [3:0]     OE_DATA_30_const_net_1;
wire   [3:0]     OE_DATA_31_const_net_1;
wire   [3:0]     OE_DATA_32_const_net_1;
wire   [3:0]     OE_DATA_33_const_net_1;
wire   [3:0]     OE_DATA_34_const_net_1;
wire   [3:0]     OE_DATA_35_const_net_1;
wire   [3:0]     OE_DATA_36_const_net_1;
wire   [3:0]     OE_DATA_37_const_net_1;
wire   [3:0]     OE_DATA_38_const_net_1;
wire   [3:0]     OE_DATA_39_const_net_1;
wire   [3:0]     OE_DATA_40_const_net_1;
wire   [3:0]     OE_DATA_41_const_net_1;
wire   [3:0]     OE_DATA_42_const_net_1;
wire   [3:0]     OE_DATA_43_const_net_1;
wire   [3:0]     OE_DATA_44_const_net_1;
wire   [3:0]     OE_DATA_45_const_net_1;
wire   [3:0]     OE_DATA_46_const_net_1;
wire   [3:0]     OE_DATA_47_const_net_1;
wire   [3:0]     OE_DATA_48_const_net_1;
wire   [3:0]     OE_DATA_49_const_net_1;
wire   [3:0]     OE_DATA_50_const_net_1;
wire   [3:0]     OE_DATA_51_const_net_1;
wire   [3:0]     OE_DATA_52_const_net_1;
wire   [3:0]     OE_DATA_53_const_net_1;
wire   [3:0]     OE_DATA_54_const_net_1;
wire   [3:0]     OE_DATA_55_const_net_1;
wire   [3:0]     OE_DATA_56_const_net_1;
wire   [3:0]     OE_DATA_57_const_net_1;
wire   [3:0]     OE_DATA_58_const_net_1;
wire   [3:0]     OE_DATA_59_const_net_1;
wire   [3:0]     OE_DATA_60_const_net_1;
wire   [3:0]     OE_DATA_61_const_net_1;
wire   [3:0]     OE_DATA_62_const_net_1;
wire   [3:0]     OE_DATA_63_const_net_1;
wire   [3:0]     OE_DATA_64_const_net_1;
wire   [3:0]     OE_DATA_65_const_net_1;
wire   [3:0]     OE_DATA_66_const_net_1;
wire   [3:0]     OE_DATA_67_const_net_1;
wire   [3:0]     OE_DATA_68_const_net_1;
wire   [3:0]     OE_DATA_69_const_net_1;
wire   [3:0]     OE_DATA_70_const_net_1;
wire   [3:0]     OE_DATA_71_const_net_1;
wire   [3:0]     OE_DATA_72_const_net_1;
wire   [3:0]     OE_DATA_73_const_net_1;
wire   [3:0]     OE_DATA_74_const_net_1;
wire   [3:0]     OE_DATA_75_const_net_1;
wire   [3:0]     OE_DATA_76_const_net_1;
wire   [3:0]     OE_DATA_77_const_net_1;
wire   [3:0]     OE_DATA_78_const_net_1;
wire   [3:0]     OE_DATA_79_const_net_1;
wire   [3:0]     OE_DATA_80_const_net_1;
wire   [3:0]     OE_DATA_81_const_net_1;
wire   [3:0]     OE_DATA_82_const_net_1;
wire   [3:0]     OE_DATA_83_const_net_1;
wire   [3:0]     OE_DATA_84_const_net_1;
wire   [3:0]     OE_DATA_85_const_net_1;
wire   [3:0]     OE_DATA_86_const_net_1;
wire   [3:0]     OE_DATA_87_const_net_1;
wire   [3:0]     OE_DATA_88_const_net_1;
wire   [3:0]     OE_DATA_89_const_net_1;
wire   [3:0]     OE_DATA_90_const_net_1;
wire   [3:0]     OE_DATA_91_const_net_1;
wire   [3:0]     OE_DATA_92_const_net_1;
wire   [3:0]     OE_DATA_93_const_net_1;
wire   [3:0]     OE_DATA_94_const_net_1;
wire   [3:0]     OE_DATA_95_const_net_1;
wire   [3:0]     OE_DATA_96_const_net_1;
wire   [3:0]     OE_DATA_97_const_net_1;
wire   [3:0]     OE_DATA_98_const_net_1;
wire   [3:0]     OE_DATA_99_const_net_1;
wire   [3:0]     OE_DATA_100_const_net_1;
wire   [3:0]     OE_DATA_101_const_net_1;
wire   [3:0]     OE_DATA_102_const_net_1;
wire   [3:0]     OE_DATA_103_const_net_1;
wire   [3:0]     OE_DATA_104_const_net_1;
wire   [3:0]     OE_DATA_105_const_net_1;
wire   [3:0]     OE_DATA_106_const_net_1;
wire   [3:0]     OE_DATA_107_const_net_1;
wire   [3:0]     OE_DATA_108_const_net_1;
wire   [3:0]     OE_DATA_109_const_net_1;
wire   [3:0]     OE_DATA_110_const_net_1;
wire   [3:0]     OE_DATA_111_const_net_1;
wire   [3:0]     OE_DATA_112_const_net_1;
wire   [3:0]     OE_DATA_113_const_net_1;
wire   [3:0]     OE_DATA_114_const_net_1;
wire   [3:0]     OE_DATA_115_const_net_1;
wire   [3:0]     OE_DATA_116_const_net_1;
wire   [3:0]     OE_DATA_117_const_net_1;
wire   [3:0]     OE_DATA_118_const_net_1;
wire   [3:0]     OE_DATA_119_const_net_1;
wire   [3:0]     OE_DATA_120_const_net_1;
wire   [3:0]     OE_DATA_121_const_net_1;
wire   [3:0]     OE_DATA_122_const_net_1;
wire   [3:0]     OE_DATA_123_const_net_1;
wire   [3:0]     OE_DATA_124_const_net_1;
wire   [3:0]     OE_DATA_125_const_net_1;
wire   [3:0]     OE_DATA_126_const_net_1;
wire   [3:0]     OE_DATA_127_const_net_1;
wire   [1:0]     RX_DQS_90_const_net_2;
wire   [2:0]     FIFO_WR_PTR_const_net_2;
wire   [2:0]     FIFO_RD_PTR_const_net_2;
wire   [2:0]     EYE_MONITOR_LANE_WIDTH_const_net_2;
wire   [3:0]     TX_DATA_1_const_net_1;
wire   [3:0]     TX_DATA_2_const_net_1;
wire   [3:0]     TX_DATA_3_const_net_1;
wire   [3:0]     TX_DATA_4_const_net_1;
wire   [3:0]     TX_DATA_5_const_net_1;
wire   [3:0]     TX_DATA_6_const_net_1;
wire   [3:0]     TX_DATA_7_const_net_1;
wire   [3:0]     TX_DATA_8_const_net_1;
wire   [3:0]     TX_DATA_9_const_net_1;
wire   [3:0]     TX_DATA_10_const_net_1;
wire   [3:0]     TX_DATA_11_const_net_1;
wire   [3:0]     TX_DATA_12_const_net_2;
wire   [3:0]     TX_DATA_13_const_net_2;
wire   [3:0]     TX_DATA_14_const_net_2;
wire   [3:0]     TX_DATA_15_const_net_2;
wire   [3:0]     TX_DATA_16_const_net_2;
wire   [3:0]     TX_DATA_17_const_net_2;
wire   [3:0]     TX_DATA_18_const_net_2;
wire   [3:0]     TX_DATA_19_const_net_2;
wire   [3:0]     TX_DATA_20_const_net_2;
wire   [3:0]     TX_DATA_21_const_net_2;
wire   [3:0]     TX_DATA_22_const_net_2;
wire   [3:0]     TX_DATA_23_const_net_2;
wire   [3:0]     TX_DATA_24_const_net_2;
wire   [3:0]     TX_DATA_25_const_net_2;
wire   [3:0]     TX_DATA_26_const_net_2;
wire   [3:0]     TX_DATA_27_const_net_2;
wire   [3:0]     TX_DATA_28_const_net_2;
wire   [3:0]     TX_DATA_29_const_net_2;
wire   [3:0]     TX_DATA_30_const_net_2;
wire   [3:0]     TX_DATA_31_const_net_2;
wire   [3:0]     TX_DATA_32_const_net_2;
wire   [3:0]     TX_DATA_33_const_net_2;
wire   [3:0]     TX_DATA_34_const_net_2;
wire   [3:0]     TX_DATA_35_const_net_2;
wire   [3:0]     TX_DATA_36_const_net_2;
wire   [3:0]     TX_DATA_37_const_net_2;
wire   [3:0]     TX_DATA_38_const_net_2;
wire   [3:0]     TX_DATA_39_const_net_2;
wire   [3:0]     TX_DATA_40_const_net_2;
wire   [3:0]     TX_DATA_41_const_net_2;
wire   [3:0]     TX_DATA_42_const_net_2;
wire   [3:0]     TX_DATA_43_const_net_2;
wire   [3:0]     TX_DATA_44_const_net_2;
wire   [3:0]     TX_DATA_45_const_net_2;
wire   [3:0]     TX_DATA_46_const_net_2;
wire   [3:0]     TX_DATA_47_const_net_2;
wire   [3:0]     TX_DATA_48_const_net_2;
wire   [3:0]     TX_DATA_49_const_net_2;
wire   [3:0]     TX_DATA_50_const_net_2;
wire   [3:0]     TX_DATA_51_const_net_2;
wire   [3:0]     TX_DATA_52_const_net_2;
wire   [3:0]     TX_DATA_53_const_net_2;
wire   [3:0]     TX_DATA_54_const_net_2;
wire   [3:0]     TX_DATA_55_const_net_2;
wire   [3:0]     TX_DATA_56_const_net_2;
wire   [3:0]     TX_DATA_57_const_net_2;
wire   [3:0]     TX_DATA_58_const_net_2;
wire   [3:0]     TX_DATA_59_const_net_2;
wire   [3:0]     TX_DATA_60_const_net_2;
wire   [3:0]     TX_DATA_61_const_net_2;
wire   [3:0]     TX_DATA_62_const_net_2;
wire   [3:0]     TX_DATA_63_const_net_2;
wire   [3:0]     TX_DATA_64_const_net_2;
wire   [3:0]     TX_DATA_65_const_net_2;
wire   [3:0]     TX_DATA_66_const_net_2;
wire   [3:0]     TX_DATA_67_const_net_2;
wire   [3:0]     TX_DATA_68_const_net_2;
wire   [3:0]     TX_DATA_69_const_net_2;
wire   [3:0]     TX_DATA_70_const_net_2;
wire   [3:0]     TX_DATA_71_const_net_2;
wire   [3:0]     TX_DATA_72_const_net_2;
wire   [3:0]     TX_DATA_73_const_net_2;
wire   [3:0]     TX_DATA_74_const_net_2;
wire   [3:0]     TX_DATA_75_const_net_2;
wire   [3:0]     TX_DATA_76_const_net_2;
wire   [3:0]     TX_DATA_77_const_net_2;
wire   [3:0]     TX_DATA_78_const_net_2;
wire   [3:0]     TX_DATA_79_const_net_2;
wire   [3:0]     TX_DATA_80_const_net_2;
wire   [3:0]     TX_DATA_81_const_net_2;
wire   [3:0]     TX_DATA_82_const_net_2;
wire   [3:0]     TX_DATA_83_const_net_2;
wire   [3:0]     TX_DATA_84_const_net_2;
wire   [3:0]     TX_DATA_85_const_net_2;
wire   [3:0]     TX_DATA_86_const_net_2;
wire   [3:0]     TX_DATA_87_const_net_2;
wire   [3:0]     TX_DATA_88_const_net_2;
wire   [3:0]     TX_DATA_89_const_net_2;
wire   [3:0]     TX_DATA_90_const_net_2;
wire   [3:0]     TX_DATA_91_const_net_2;
wire   [3:0]     TX_DATA_92_const_net_2;
wire   [3:0]     TX_DATA_93_const_net_2;
wire   [3:0]     TX_DATA_94_const_net_2;
wire   [3:0]     TX_DATA_95_const_net_2;
wire   [3:0]     TX_DATA_96_const_net_2;
wire   [3:0]     TX_DATA_97_const_net_2;
wire   [3:0]     TX_DATA_98_const_net_2;
wire   [3:0]     TX_DATA_99_const_net_2;
wire   [3:0]     TX_DATA_100_const_net_2;
wire   [3:0]     TX_DATA_101_const_net_2;
wire   [3:0]     TX_DATA_102_const_net_2;
wire   [3:0]     TX_DATA_103_const_net_2;
wire   [3:0]     TX_DATA_104_const_net_2;
wire   [3:0]     TX_DATA_105_const_net_2;
wire   [3:0]     TX_DATA_106_const_net_2;
wire   [3:0]     TX_DATA_107_const_net_2;
wire   [3:0]     TX_DATA_108_const_net_2;
wire   [3:0]     TX_DATA_109_const_net_2;
wire   [3:0]     TX_DATA_110_const_net_2;
wire   [3:0]     TX_DATA_111_const_net_2;
wire   [3:0]     TX_DATA_112_const_net_2;
wire   [3:0]     TX_DATA_113_const_net_2;
wire   [3:0]     TX_DATA_114_const_net_2;
wire   [3:0]     TX_DATA_115_const_net_2;
wire   [3:0]     TX_DATA_116_const_net_2;
wire   [3:0]     TX_DATA_117_const_net_2;
wire   [3:0]     TX_DATA_118_const_net_2;
wire   [3:0]     TX_DATA_119_const_net_2;
wire   [3:0]     TX_DATA_120_const_net_2;
wire   [3:0]     TX_DATA_121_const_net_2;
wire   [3:0]     TX_DATA_122_const_net_2;
wire   [3:0]     TX_DATA_123_const_net_2;
wire   [3:0]     TX_DATA_124_const_net_2;
wire   [3:0]     TX_DATA_125_const_net_2;
wire   [3:0]     TX_DATA_126_const_net_2;
wire   [3:0]     TX_DATA_127_const_net_2;
wire   [3:0]     OE_DATA_1_const_net_4;
wire   [3:0]     OE_DATA_2_const_net_2;
wire   [3:0]     OE_DATA_3_const_net_2;
wire   [3:0]     OE_DATA_4_const_net_2;
wire   [3:0]     OE_DATA_5_const_net_2;
wire   [3:0]     OE_DATA_6_const_net_2;
wire   [3:0]     OE_DATA_7_const_net_2;
wire   [3:0]     OE_DATA_8_const_net_2;
wire   [3:0]     OE_DATA_9_const_net_2;
wire   [3:0]     OE_DATA_10_const_net_2;
wire   [3:0]     OE_DATA_11_const_net_2;
wire   [3:0]     OE_DATA_12_const_net_2;
wire   [3:0]     OE_DATA_13_const_net_2;
wire   [3:0]     OE_DATA_14_const_net_2;
wire   [3:0]     OE_DATA_15_const_net_2;
wire   [3:0]     OE_DATA_16_const_net_2;
wire   [3:0]     OE_DATA_17_const_net_2;
wire   [3:0]     OE_DATA_18_const_net_2;
wire   [3:0]     OE_DATA_19_const_net_2;
wire   [3:0]     OE_DATA_20_const_net_2;
wire   [3:0]     OE_DATA_21_const_net_2;
wire   [3:0]     OE_DATA_22_const_net_2;
wire   [3:0]     OE_DATA_23_const_net_2;
wire   [3:0]     OE_DATA_24_const_net_2;
wire   [3:0]     OE_DATA_25_const_net_2;
wire   [3:0]     OE_DATA_26_const_net_2;
wire   [3:0]     OE_DATA_27_const_net_2;
wire   [3:0]     OE_DATA_28_const_net_2;
wire   [3:0]     OE_DATA_29_const_net_2;
wire   [3:0]     OE_DATA_30_const_net_2;
wire   [3:0]     OE_DATA_31_const_net_2;
wire   [3:0]     OE_DATA_32_const_net_2;
wire   [3:0]     OE_DATA_33_const_net_2;
wire   [3:0]     OE_DATA_34_const_net_2;
wire   [3:0]     OE_DATA_35_const_net_2;
wire   [3:0]     OE_DATA_36_const_net_2;
wire   [3:0]     OE_DATA_37_const_net_2;
wire   [3:0]     OE_DATA_38_const_net_2;
wire   [3:0]     OE_DATA_39_const_net_2;
wire   [3:0]     OE_DATA_40_const_net_2;
wire   [3:0]     OE_DATA_41_const_net_2;
wire   [3:0]     OE_DATA_42_const_net_2;
wire   [3:0]     OE_DATA_43_const_net_2;
wire   [3:0]     OE_DATA_44_const_net_2;
wire   [3:0]     OE_DATA_45_const_net_2;
wire   [3:0]     OE_DATA_46_const_net_2;
wire   [3:0]     OE_DATA_47_const_net_2;
wire   [3:0]     OE_DATA_48_const_net_2;
wire   [3:0]     OE_DATA_49_const_net_2;
wire   [3:0]     OE_DATA_50_const_net_2;
wire   [3:0]     OE_DATA_51_const_net_2;
wire   [3:0]     OE_DATA_52_const_net_2;
wire   [3:0]     OE_DATA_53_const_net_2;
wire   [3:0]     OE_DATA_54_const_net_2;
wire   [3:0]     OE_DATA_55_const_net_2;
wire   [3:0]     OE_DATA_56_const_net_2;
wire   [3:0]     OE_DATA_57_const_net_2;
wire   [3:0]     OE_DATA_58_const_net_2;
wire   [3:0]     OE_DATA_59_const_net_2;
wire   [3:0]     OE_DATA_60_const_net_2;
wire   [3:0]     OE_DATA_61_const_net_2;
wire   [3:0]     OE_DATA_62_const_net_2;
wire   [3:0]     OE_DATA_63_const_net_2;
wire   [3:0]     OE_DATA_64_const_net_2;
wire   [3:0]     OE_DATA_65_const_net_2;
wire   [3:0]     OE_DATA_66_const_net_2;
wire   [3:0]     OE_DATA_67_const_net_2;
wire   [3:0]     OE_DATA_68_const_net_2;
wire   [3:0]     OE_DATA_69_const_net_2;
wire   [3:0]     OE_DATA_70_const_net_2;
wire   [3:0]     OE_DATA_71_const_net_2;
wire   [3:0]     OE_DATA_72_const_net_2;
wire   [3:0]     OE_DATA_73_const_net_2;
wire   [3:0]     OE_DATA_74_const_net_2;
wire   [3:0]     OE_DATA_75_const_net_2;
wire   [3:0]     OE_DATA_76_const_net_2;
wire   [3:0]     OE_DATA_77_const_net_2;
wire   [3:0]     OE_DATA_78_const_net_2;
wire   [3:0]     OE_DATA_79_const_net_2;
wire   [3:0]     OE_DATA_80_const_net_2;
wire   [3:0]     OE_DATA_81_const_net_2;
wire   [3:0]     OE_DATA_82_const_net_2;
wire   [3:0]     OE_DATA_83_const_net_2;
wire   [3:0]     OE_DATA_84_const_net_2;
wire   [3:0]     OE_DATA_85_const_net_2;
wire   [3:0]     OE_DATA_86_const_net_2;
wire   [3:0]     OE_DATA_87_const_net_2;
wire   [3:0]     OE_DATA_88_const_net_2;
wire   [3:0]     OE_DATA_89_const_net_2;
wire   [3:0]     OE_DATA_90_const_net_2;
wire   [3:0]     OE_DATA_91_const_net_2;
wire   [3:0]     OE_DATA_92_const_net_2;
wire   [3:0]     OE_DATA_93_const_net_2;
wire   [3:0]     OE_DATA_94_const_net_2;
wire   [3:0]     OE_DATA_95_const_net_2;
wire   [3:0]     OE_DATA_96_const_net_2;
wire   [3:0]     OE_DATA_97_const_net_2;
wire   [3:0]     OE_DATA_98_const_net_2;
wire   [3:0]     OE_DATA_99_const_net_2;
wire   [3:0]     OE_DATA_100_const_net_2;
wire   [3:0]     OE_DATA_101_const_net_2;
wire   [3:0]     OE_DATA_102_const_net_2;
wire   [3:0]     OE_DATA_103_const_net_2;
wire   [3:0]     OE_DATA_104_const_net_2;
wire   [3:0]     OE_DATA_105_const_net_2;
wire   [3:0]     OE_DATA_106_const_net_2;
wire   [3:0]     OE_DATA_107_const_net_2;
wire   [3:0]     OE_DATA_108_const_net_2;
wire   [3:0]     OE_DATA_109_const_net_2;
wire   [3:0]     OE_DATA_110_const_net_2;
wire   [3:0]     OE_DATA_111_const_net_2;
wire   [3:0]     OE_DATA_112_const_net_2;
wire   [3:0]     OE_DATA_113_const_net_2;
wire   [3:0]     OE_DATA_114_const_net_2;
wire   [3:0]     OE_DATA_115_const_net_2;
wire   [3:0]     OE_DATA_116_const_net_2;
wire   [3:0]     OE_DATA_117_const_net_2;
wire   [3:0]     OE_DATA_118_const_net_2;
wire   [3:0]     OE_DATA_119_const_net_2;
wire   [3:0]     OE_DATA_120_const_net_2;
wire   [3:0]     OE_DATA_121_const_net_2;
wire   [3:0]     OE_DATA_122_const_net_2;
wire   [3:0]     OE_DATA_123_const_net_2;
wire   [3:0]     OE_DATA_124_const_net_2;
wire   [3:0]     OE_DATA_125_const_net_2;
wire   [3:0]     OE_DATA_126_const_net_2;
wire   [3:0]     OE_DATA_127_const_net_2;
wire   [1:0]     RX_DQS_90_const_net_3;
wire   [2:0]     FIFO_WR_PTR_const_net_3;
wire   [2:0]     FIFO_RD_PTR_const_net_3;
wire   [2:0]     EYE_MONITOR_LANE_WIDTH_const_net_3;
wire   [3:0]     TX_DATA_1_const_net_2;
wire   [3:0]     TX_DATA_2_const_net_2;
wire   [3:0]     TX_DATA_3_const_net_2;
wire   [3:0]     TX_DATA_4_const_net_2;
wire   [3:0]     TX_DATA_5_const_net_2;
wire   [3:0]     TX_DATA_6_const_net_2;
wire   [3:0]     TX_DATA_7_const_net_2;
wire   [3:0]     TX_DATA_8_const_net_2;
wire   [3:0]     TX_DATA_9_const_net_2;
wire   [3:0]     TX_DATA_10_const_net_2;
wire   [3:0]     TX_DATA_11_const_net_2;
wire   [3:0]     TX_DATA_12_const_net_3;
wire   [3:0]     TX_DATA_13_const_net_3;
wire   [3:0]     TX_DATA_14_const_net_3;
wire   [3:0]     TX_DATA_15_const_net_3;
wire   [3:0]     TX_DATA_16_const_net_3;
wire   [3:0]     TX_DATA_17_const_net_3;
wire   [3:0]     TX_DATA_18_const_net_3;
wire   [3:0]     TX_DATA_19_const_net_3;
wire   [3:0]     TX_DATA_20_const_net_3;
wire   [3:0]     TX_DATA_21_const_net_3;
wire   [3:0]     TX_DATA_22_const_net_3;
wire   [3:0]     TX_DATA_23_const_net_3;
wire   [3:0]     TX_DATA_24_const_net_3;
wire   [3:0]     TX_DATA_25_const_net_3;
wire   [3:0]     TX_DATA_26_const_net_3;
wire   [3:0]     TX_DATA_27_const_net_3;
wire   [3:0]     TX_DATA_28_const_net_3;
wire   [3:0]     TX_DATA_29_const_net_3;
wire   [3:0]     TX_DATA_30_const_net_3;
wire   [3:0]     TX_DATA_31_const_net_3;
wire   [3:0]     TX_DATA_32_const_net_3;
wire   [3:0]     TX_DATA_33_const_net_3;
wire   [3:0]     TX_DATA_34_const_net_3;
wire   [3:0]     TX_DATA_35_const_net_3;
wire   [3:0]     TX_DATA_36_const_net_3;
wire   [3:0]     TX_DATA_37_const_net_3;
wire   [3:0]     TX_DATA_38_const_net_3;
wire   [3:0]     TX_DATA_39_const_net_3;
wire   [3:0]     TX_DATA_40_const_net_3;
wire   [3:0]     TX_DATA_41_const_net_3;
wire   [3:0]     TX_DATA_42_const_net_3;
wire   [3:0]     TX_DATA_43_const_net_3;
wire   [3:0]     TX_DATA_44_const_net_3;
wire   [3:0]     TX_DATA_45_const_net_3;
wire   [3:0]     TX_DATA_46_const_net_3;
wire   [3:0]     TX_DATA_47_const_net_3;
wire   [3:0]     TX_DATA_48_const_net_3;
wire   [3:0]     TX_DATA_49_const_net_3;
wire   [3:0]     TX_DATA_50_const_net_3;
wire   [3:0]     TX_DATA_51_const_net_3;
wire   [3:0]     TX_DATA_52_const_net_3;
wire   [3:0]     TX_DATA_53_const_net_3;
wire   [3:0]     TX_DATA_54_const_net_3;
wire   [3:0]     TX_DATA_55_const_net_3;
wire   [3:0]     TX_DATA_56_const_net_3;
wire   [3:0]     TX_DATA_57_const_net_3;
wire   [3:0]     TX_DATA_58_const_net_3;
wire   [3:0]     TX_DATA_59_const_net_3;
wire   [3:0]     TX_DATA_60_const_net_3;
wire   [3:0]     TX_DATA_61_const_net_3;
wire   [3:0]     TX_DATA_62_const_net_3;
wire   [3:0]     TX_DATA_63_const_net_3;
wire   [3:0]     TX_DATA_64_const_net_3;
wire   [3:0]     TX_DATA_65_const_net_3;
wire   [3:0]     TX_DATA_66_const_net_3;
wire   [3:0]     TX_DATA_67_const_net_3;
wire   [3:0]     TX_DATA_68_const_net_3;
wire   [3:0]     TX_DATA_69_const_net_3;
wire   [3:0]     TX_DATA_70_const_net_3;
wire   [3:0]     TX_DATA_71_const_net_3;
wire   [3:0]     TX_DATA_72_const_net_3;
wire   [3:0]     TX_DATA_73_const_net_3;
wire   [3:0]     TX_DATA_74_const_net_3;
wire   [3:0]     TX_DATA_75_const_net_3;
wire   [3:0]     TX_DATA_76_const_net_3;
wire   [3:0]     TX_DATA_77_const_net_3;
wire   [3:0]     TX_DATA_78_const_net_3;
wire   [3:0]     TX_DATA_79_const_net_3;
wire   [3:0]     TX_DATA_80_const_net_3;
wire   [3:0]     TX_DATA_81_const_net_3;
wire   [3:0]     TX_DATA_82_const_net_3;
wire   [3:0]     TX_DATA_83_const_net_3;
wire   [3:0]     TX_DATA_84_const_net_3;
wire   [3:0]     TX_DATA_85_const_net_3;
wire   [3:0]     TX_DATA_86_const_net_3;
wire   [3:0]     TX_DATA_87_const_net_3;
wire   [3:0]     TX_DATA_88_const_net_3;
wire   [3:0]     TX_DATA_89_const_net_3;
wire   [3:0]     TX_DATA_90_const_net_3;
wire   [3:0]     TX_DATA_91_const_net_3;
wire   [3:0]     TX_DATA_92_const_net_3;
wire   [3:0]     TX_DATA_93_const_net_3;
wire   [3:0]     TX_DATA_94_const_net_3;
wire   [3:0]     TX_DATA_95_const_net_3;
wire   [3:0]     TX_DATA_96_const_net_3;
wire   [3:0]     TX_DATA_97_const_net_3;
wire   [3:0]     TX_DATA_98_const_net_3;
wire   [3:0]     TX_DATA_99_const_net_3;
wire   [3:0]     TX_DATA_100_const_net_3;
wire   [3:0]     TX_DATA_101_const_net_3;
wire   [3:0]     TX_DATA_102_const_net_3;
wire   [3:0]     TX_DATA_103_const_net_3;
wire   [3:0]     TX_DATA_104_const_net_3;
wire   [3:0]     TX_DATA_105_const_net_3;
wire   [3:0]     TX_DATA_106_const_net_3;
wire   [3:0]     TX_DATA_107_const_net_3;
wire   [3:0]     TX_DATA_108_const_net_3;
wire   [3:0]     TX_DATA_109_const_net_3;
wire   [3:0]     TX_DATA_110_const_net_3;
wire   [3:0]     TX_DATA_111_const_net_3;
wire   [3:0]     TX_DATA_112_const_net_3;
wire   [3:0]     TX_DATA_113_const_net_3;
wire   [3:0]     TX_DATA_114_const_net_3;
wire   [3:0]     TX_DATA_115_const_net_3;
wire   [3:0]     TX_DATA_116_const_net_3;
wire   [3:0]     TX_DATA_117_const_net_3;
wire   [3:0]     TX_DATA_118_const_net_3;
wire   [3:0]     TX_DATA_119_const_net_3;
wire   [3:0]     TX_DATA_120_const_net_3;
wire   [3:0]     TX_DATA_121_const_net_3;
wire   [3:0]     TX_DATA_122_const_net_3;
wire   [3:0]     TX_DATA_123_const_net_3;
wire   [3:0]     TX_DATA_124_const_net_3;
wire   [3:0]     TX_DATA_125_const_net_3;
wire   [3:0]     TX_DATA_126_const_net_3;
wire   [3:0]     TX_DATA_127_const_net_3;
wire   [3:0]     OE_DATA_1_const_net_5;
wire   [3:0]     OE_DATA_2_const_net_3;
wire   [3:0]     OE_DATA_3_const_net_3;
wire   [3:0]     OE_DATA_4_const_net_3;
wire   [3:0]     OE_DATA_5_const_net_3;
wire   [3:0]     OE_DATA_6_const_net_3;
wire   [3:0]     OE_DATA_7_const_net_3;
wire   [3:0]     OE_DATA_8_const_net_3;
wire   [3:0]     OE_DATA_9_const_net_3;
wire   [3:0]     OE_DATA_10_const_net_3;
wire   [3:0]     OE_DATA_11_const_net_3;
wire   [3:0]     OE_DATA_12_const_net_3;
wire   [3:0]     OE_DATA_13_const_net_3;
wire   [3:0]     OE_DATA_14_const_net_3;
wire   [3:0]     OE_DATA_15_const_net_3;
wire   [3:0]     OE_DATA_16_const_net_3;
wire   [3:0]     OE_DATA_17_const_net_3;
wire   [3:0]     OE_DATA_18_const_net_3;
wire   [3:0]     OE_DATA_19_const_net_3;
wire   [3:0]     OE_DATA_20_const_net_3;
wire   [3:0]     OE_DATA_21_const_net_3;
wire   [3:0]     OE_DATA_22_const_net_3;
wire   [3:0]     OE_DATA_23_const_net_3;
wire   [3:0]     OE_DATA_24_const_net_3;
wire   [3:0]     OE_DATA_25_const_net_3;
wire   [3:0]     OE_DATA_26_const_net_3;
wire   [3:0]     OE_DATA_27_const_net_3;
wire   [3:0]     OE_DATA_28_const_net_3;
wire   [3:0]     OE_DATA_29_const_net_3;
wire   [3:0]     OE_DATA_30_const_net_3;
wire   [3:0]     OE_DATA_31_const_net_3;
wire   [3:0]     OE_DATA_32_const_net_3;
wire   [3:0]     OE_DATA_33_const_net_3;
wire   [3:0]     OE_DATA_34_const_net_3;
wire   [3:0]     OE_DATA_35_const_net_3;
wire   [3:0]     OE_DATA_36_const_net_3;
wire   [3:0]     OE_DATA_37_const_net_3;
wire   [3:0]     OE_DATA_38_const_net_3;
wire   [3:0]     OE_DATA_39_const_net_3;
wire   [3:0]     OE_DATA_40_const_net_3;
wire   [3:0]     OE_DATA_41_const_net_3;
wire   [3:0]     OE_DATA_42_const_net_3;
wire   [3:0]     OE_DATA_43_const_net_3;
wire   [3:0]     OE_DATA_44_const_net_3;
wire   [3:0]     OE_DATA_45_const_net_3;
wire   [3:0]     OE_DATA_46_const_net_3;
wire   [3:0]     OE_DATA_47_const_net_3;
wire   [3:0]     OE_DATA_48_const_net_3;
wire   [3:0]     OE_DATA_49_const_net_3;
wire   [3:0]     OE_DATA_50_const_net_3;
wire   [3:0]     OE_DATA_51_const_net_3;
wire   [3:0]     OE_DATA_52_const_net_3;
wire   [3:0]     OE_DATA_53_const_net_3;
wire   [3:0]     OE_DATA_54_const_net_3;
wire   [3:0]     OE_DATA_55_const_net_3;
wire   [3:0]     OE_DATA_56_const_net_3;
wire   [3:0]     OE_DATA_57_const_net_3;
wire   [3:0]     OE_DATA_58_const_net_3;
wire   [3:0]     OE_DATA_59_const_net_3;
wire   [3:0]     OE_DATA_60_const_net_3;
wire   [3:0]     OE_DATA_61_const_net_3;
wire   [3:0]     OE_DATA_62_const_net_3;
wire   [3:0]     OE_DATA_63_const_net_3;
wire   [3:0]     OE_DATA_64_const_net_3;
wire   [3:0]     OE_DATA_65_const_net_3;
wire   [3:0]     OE_DATA_66_const_net_3;
wire   [3:0]     OE_DATA_67_const_net_3;
wire   [3:0]     OE_DATA_68_const_net_3;
wire   [3:0]     OE_DATA_69_const_net_3;
wire   [3:0]     OE_DATA_70_const_net_3;
wire   [3:0]     OE_DATA_71_const_net_3;
wire   [3:0]     OE_DATA_72_const_net_3;
wire   [3:0]     OE_DATA_73_const_net_3;
wire   [3:0]     OE_DATA_74_const_net_3;
wire   [3:0]     OE_DATA_75_const_net_3;
wire   [3:0]     OE_DATA_76_const_net_3;
wire   [3:0]     OE_DATA_77_const_net_3;
wire   [3:0]     OE_DATA_78_const_net_3;
wire   [3:0]     OE_DATA_79_const_net_3;
wire   [3:0]     OE_DATA_80_const_net_3;
wire   [3:0]     OE_DATA_81_const_net_3;
wire   [3:0]     OE_DATA_82_const_net_3;
wire   [3:0]     OE_DATA_83_const_net_3;
wire   [3:0]     OE_DATA_84_const_net_3;
wire   [3:0]     OE_DATA_85_const_net_3;
wire   [3:0]     OE_DATA_86_const_net_3;
wire   [3:0]     OE_DATA_87_const_net_3;
wire   [3:0]     OE_DATA_88_const_net_3;
wire   [3:0]     OE_DATA_89_const_net_3;
wire   [3:0]     OE_DATA_90_const_net_3;
wire   [3:0]     OE_DATA_91_const_net_3;
wire   [3:0]     OE_DATA_92_const_net_3;
wire   [3:0]     OE_DATA_93_const_net_3;
wire   [3:0]     OE_DATA_94_const_net_3;
wire   [3:0]     OE_DATA_95_const_net_3;
wire   [3:0]     OE_DATA_96_const_net_3;
wire   [3:0]     OE_DATA_97_const_net_3;
wire   [3:0]     OE_DATA_98_const_net_3;
wire   [3:0]     OE_DATA_99_const_net_3;
wire   [3:0]     OE_DATA_100_const_net_3;
wire   [3:0]     OE_DATA_101_const_net_3;
wire   [3:0]     OE_DATA_102_const_net_3;
wire   [3:0]     OE_DATA_103_const_net_3;
wire   [3:0]     OE_DATA_104_const_net_3;
wire   [3:0]     OE_DATA_105_const_net_3;
wire   [3:0]     OE_DATA_106_const_net_3;
wire   [3:0]     OE_DATA_107_const_net_3;
wire   [3:0]     OE_DATA_108_const_net_3;
wire   [3:0]     OE_DATA_109_const_net_3;
wire   [3:0]     OE_DATA_110_const_net_3;
wire   [3:0]     OE_DATA_111_const_net_3;
wire   [3:0]     OE_DATA_112_const_net_3;
wire   [3:0]     OE_DATA_113_const_net_3;
wire   [3:0]     OE_DATA_114_const_net_3;
wire   [3:0]     OE_DATA_115_const_net_3;
wire   [3:0]     OE_DATA_116_const_net_3;
wire   [3:0]     OE_DATA_117_const_net_3;
wire   [3:0]     OE_DATA_118_const_net_3;
wire   [3:0]     OE_DATA_119_const_net_3;
wire   [3:0]     OE_DATA_120_const_net_3;
wire   [3:0]     OE_DATA_121_const_net_3;
wire   [3:0]     OE_DATA_122_const_net_3;
wire   [3:0]     OE_DATA_123_const_net_3;
wire   [3:0]     OE_DATA_124_const_net_3;
wire   [3:0]     OE_DATA_125_const_net_3;
wire   [3:0]     OE_DATA_126_const_net_3;
wire   [3:0]     OE_DATA_127_const_net_3;
wire   [1:0]     RX_DQS_90_const_net_4;
wire   [2:0]     FIFO_WR_PTR_const_net_4;
wire   [2:0]     FIFO_RD_PTR_const_net_4;
wire   [2:0]     EYE_MONITOR_LANE_WIDTH_const_net_4;
wire   [3:0]     TX_DATA_2_const_net_3;
wire   [3:0]     TX_DATA_3_const_net_3;
wire   [3:0]     TX_DATA_4_const_net_3;
wire   [3:0]     TX_DATA_5_const_net_3;
wire   [3:0]     TX_DATA_6_const_net_3;
wire   [3:0]     TX_DATA_7_const_net_3;
wire   [3:0]     TX_DATA_8_const_net_3;
wire   [3:0]     TX_DATA_9_const_net_3;
wire   [3:0]     TX_DATA_10_const_net_3;
wire   [3:0]     TX_DATA_11_const_net_3;
wire   [3:0]     TX_DATA_12_const_net_4;
wire   [3:0]     TX_DATA_13_const_net_4;
wire   [3:0]     TX_DATA_14_const_net_4;
wire   [3:0]     TX_DATA_15_const_net_4;
wire   [3:0]     TX_DATA_16_const_net_4;
wire   [3:0]     TX_DATA_17_const_net_4;
wire   [3:0]     TX_DATA_18_const_net_4;
wire   [3:0]     TX_DATA_19_const_net_4;
wire   [3:0]     TX_DATA_20_const_net_4;
wire   [3:0]     TX_DATA_21_const_net_4;
wire   [3:0]     TX_DATA_22_const_net_4;
wire   [3:0]     TX_DATA_23_const_net_4;
wire   [3:0]     TX_DATA_24_const_net_4;
wire   [3:0]     TX_DATA_25_const_net_4;
wire   [3:0]     TX_DATA_26_const_net_4;
wire   [3:0]     TX_DATA_27_const_net_4;
wire   [3:0]     TX_DATA_28_const_net_4;
wire   [3:0]     TX_DATA_29_const_net_4;
wire   [3:0]     TX_DATA_30_const_net_4;
wire   [3:0]     TX_DATA_31_const_net_4;
wire   [3:0]     TX_DATA_32_const_net_4;
wire   [3:0]     TX_DATA_33_const_net_4;
wire   [3:0]     TX_DATA_34_const_net_4;
wire   [3:0]     TX_DATA_35_const_net_4;
wire   [3:0]     TX_DATA_36_const_net_4;
wire   [3:0]     TX_DATA_37_const_net_4;
wire   [3:0]     TX_DATA_38_const_net_4;
wire   [3:0]     TX_DATA_39_const_net_4;
wire   [3:0]     TX_DATA_40_const_net_4;
wire   [3:0]     TX_DATA_41_const_net_4;
wire   [3:0]     TX_DATA_42_const_net_4;
wire   [3:0]     TX_DATA_43_const_net_4;
wire   [3:0]     TX_DATA_44_const_net_4;
wire   [3:0]     TX_DATA_45_const_net_4;
wire   [3:0]     TX_DATA_46_const_net_4;
wire   [3:0]     TX_DATA_47_const_net_4;
wire   [3:0]     TX_DATA_48_const_net_4;
wire   [3:0]     TX_DATA_49_const_net_4;
wire   [3:0]     TX_DATA_50_const_net_4;
wire   [3:0]     TX_DATA_51_const_net_4;
wire   [3:0]     TX_DATA_52_const_net_4;
wire   [3:0]     TX_DATA_53_const_net_4;
wire   [3:0]     TX_DATA_54_const_net_4;
wire   [3:0]     TX_DATA_55_const_net_4;
wire   [3:0]     TX_DATA_56_const_net_4;
wire   [3:0]     TX_DATA_57_const_net_4;
wire   [3:0]     TX_DATA_58_const_net_4;
wire   [3:0]     TX_DATA_59_const_net_4;
wire   [3:0]     TX_DATA_60_const_net_4;
wire   [3:0]     TX_DATA_61_const_net_4;
wire   [3:0]     TX_DATA_62_const_net_4;
wire   [3:0]     TX_DATA_63_const_net_4;
wire   [3:0]     TX_DATA_64_const_net_4;
wire   [3:0]     TX_DATA_65_const_net_4;
wire   [3:0]     TX_DATA_66_const_net_4;
wire   [3:0]     TX_DATA_67_const_net_4;
wire   [3:0]     TX_DATA_68_const_net_4;
wire   [3:0]     TX_DATA_69_const_net_4;
wire   [3:0]     TX_DATA_70_const_net_4;
wire   [3:0]     TX_DATA_71_const_net_4;
wire   [3:0]     TX_DATA_72_const_net_4;
wire   [3:0]     TX_DATA_73_const_net_4;
wire   [3:0]     TX_DATA_74_const_net_4;
wire   [3:0]     TX_DATA_75_const_net_4;
wire   [3:0]     TX_DATA_76_const_net_4;
wire   [3:0]     TX_DATA_77_const_net_4;
wire   [3:0]     TX_DATA_78_const_net_4;
wire   [3:0]     TX_DATA_79_const_net_4;
wire   [3:0]     TX_DATA_80_const_net_4;
wire   [3:0]     TX_DATA_81_const_net_4;
wire   [3:0]     TX_DATA_82_const_net_4;
wire   [3:0]     TX_DATA_83_const_net_4;
wire   [3:0]     TX_DATA_84_const_net_4;
wire   [3:0]     TX_DATA_85_const_net_4;
wire   [3:0]     TX_DATA_86_const_net_4;
wire   [3:0]     TX_DATA_87_const_net_4;
wire   [3:0]     TX_DATA_88_const_net_4;
wire   [3:0]     TX_DATA_89_const_net_4;
wire   [3:0]     TX_DATA_90_const_net_4;
wire   [3:0]     TX_DATA_91_const_net_4;
wire   [3:0]     TX_DATA_92_const_net_4;
wire   [3:0]     TX_DATA_93_const_net_4;
wire   [3:0]     TX_DATA_94_const_net_4;
wire   [3:0]     TX_DATA_95_const_net_4;
wire   [3:0]     TX_DATA_96_const_net_4;
wire   [3:0]     TX_DATA_97_const_net_4;
wire   [3:0]     TX_DATA_98_const_net_4;
wire   [3:0]     TX_DATA_99_const_net_4;
wire   [3:0]     TX_DATA_100_const_net_4;
wire   [3:0]     TX_DATA_101_const_net_4;
wire   [3:0]     TX_DATA_102_const_net_4;
wire   [3:0]     TX_DATA_103_const_net_4;
wire   [3:0]     TX_DATA_104_const_net_4;
wire   [3:0]     TX_DATA_105_const_net_4;
wire   [3:0]     TX_DATA_106_const_net_4;
wire   [3:0]     TX_DATA_107_const_net_4;
wire   [3:0]     TX_DATA_108_const_net_4;
wire   [3:0]     TX_DATA_109_const_net_4;
wire   [3:0]     TX_DATA_110_const_net_4;
wire   [3:0]     TX_DATA_111_const_net_4;
wire   [3:0]     TX_DATA_112_const_net_4;
wire   [3:0]     TX_DATA_113_const_net_4;
wire   [3:0]     TX_DATA_114_const_net_4;
wire   [3:0]     TX_DATA_115_const_net_4;
wire   [3:0]     TX_DATA_116_const_net_4;
wire   [3:0]     TX_DATA_117_const_net_4;
wire   [3:0]     TX_DATA_118_const_net_4;
wire   [3:0]     TX_DATA_119_const_net_4;
wire   [3:0]     TX_DATA_120_const_net_4;
wire   [3:0]     TX_DATA_121_const_net_4;
wire   [3:0]     TX_DATA_122_const_net_4;
wire   [3:0]     TX_DATA_123_const_net_4;
wire   [3:0]     TX_DATA_124_const_net_4;
wire   [3:0]     TX_DATA_125_const_net_4;
wire   [3:0]     TX_DATA_126_const_net_4;
wire   [3:0]     TX_DATA_127_const_net_4;
wire   [3:0]     OE_DATA_2_const_net_4;
wire   [3:0]     OE_DATA_3_const_net_4;
wire   [3:0]     OE_DATA_4_const_net_4;
wire   [3:0]     OE_DATA_5_const_net_4;
wire   [3:0]     OE_DATA_6_const_net_4;
wire   [3:0]     OE_DATA_7_const_net_4;
wire   [3:0]     OE_DATA_8_const_net_4;
wire   [3:0]     OE_DATA_9_const_net_4;
wire   [3:0]     OE_DATA_10_const_net_4;
wire   [3:0]     OE_DATA_11_const_net_4;
wire   [3:0]     OE_DATA_12_const_net_4;
wire   [3:0]     OE_DATA_13_const_net_4;
wire   [3:0]     OE_DATA_14_const_net_4;
wire   [3:0]     OE_DATA_15_const_net_4;
wire   [3:0]     OE_DATA_16_const_net_4;
wire   [3:0]     OE_DATA_17_const_net_4;
wire   [3:0]     OE_DATA_18_const_net_4;
wire   [3:0]     OE_DATA_19_const_net_4;
wire   [3:0]     OE_DATA_20_const_net_4;
wire   [3:0]     OE_DATA_21_const_net_4;
wire   [3:0]     OE_DATA_22_const_net_4;
wire   [3:0]     OE_DATA_23_const_net_4;
wire   [3:0]     OE_DATA_24_const_net_4;
wire   [3:0]     OE_DATA_25_const_net_4;
wire   [3:0]     OE_DATA_26_const_net_4;
wire   [3:0]     OE_DATA_27_const_net_4;
wire   [3:0]     OE_DATA_28_const_net_4;
wire   [3:0]     OE_DATA_29_const_net_4;
wire   [3:0]     OE_DATA_30_const_net_4;
wire   [3:0]     OE_DATA_31_const_net_4;
wire   [3:0]     OE_DATA_32_const_net_4;
wire   [3:0]     OE_DATA_33_const_net_4;
wire   [3:0]     OE_DATA_34_const_net_4;
wire   [3:0]     OE_DATA_35_const_net_4;
wire   [3:0]     OE_DATA_36_const_net_4;
wire   [3:0]     OE_DATA_37_const_net_4;
wire   [3:0]     OE_DATA_38_const_net_4;
wire   [3:0]     OE_DATA_39_const_net_4;
wire   [3:0]     OE_DATA_40_const_net_4;
wire   [3:0]     OE_DATA_41_const_net_4;
wire   [3:0]     OE_DATA_42_const_net_4;
wire   [3:0]     OE_DATA_43_const_net_4;
wire   [3:0]     OE_DATA_44_const_net_4;
wire   [3:0]     OE_DATA_45_const_net_4;
wire   [3:0]     OE_DATA_46_const_net_4;
wire   [3:0]     OE_DATA_47_const_net_4;
wire   [3:0]     OE_DATA_48_const_net_4;
wire   [3:0]     OE_DATA_49_const_net_4;
wire   [3:0]     OE_DATA_50_const_net_4;
wire   [3:0]     OE_DATA_51_const_net_4;
wire   [3:0]     OE_DATA_52_const_net_4;
wire   [3:0]     OE_DATA_53_const_net_4;
wire   [3:0]     OE_DATA_54_const_net_4;
wire   [3:0]     OE_DATA_55_const_net_4;
wire   [3:0]     OE_DATA_56_const_net_4;
wire   [3:0]     OE_DATA_57_const_net_4;
wire   [3:0]     OE_DATA_58_const_net_4;
wire   [3:0]     OE_DATA_59_const_net_4;
wire   [3:0]     OE_DATA_60_const_net_4;
wire   [3:0]     OE_DATA_61_const_net_4;
wire   [3:0]     OE_DATA_62_const_net_4;
wire   [3:0]     OE_DATA_63_const_net_4;
wire   [3:0]     OE_DATA_64_const_net_4;
wire   [3:0]     OE_DATA_65_const_net_4;
wire   [3:0]     OE_DATA_66_const_net_4;
wire   [3:0]     OE_DATA_67_const_net_4;
wire   [3:0]     OE_DATA_68_const_net_4;
wire   [3:0]     OE_DATA_69_const_net_4;
wire   [3:0]     OE_DATA_70_const_net_4;
wire   [3:0]     OE_DATA_71_const_net_4;
wire   [3:0]     OE_DATA_72_const_net_4;
wire   [3:0]     OE_DATA_73_const_net_4;
wire   [3:0]     OE_DATA_74_const_net_4;
wire   [3:0]     OE_DATA_75_const_net_4;
wire   [3:0]     OE_DATA_76_const_net_4;
wire   [3:0]     OE_DATA_77_const_net_4;
wire   [3:0]     OE_DATA_78_const_net_4;
wire   [3:0]     OE_DATA_79_const_net_4;
wire   [3:0]     OE_DATA_80_const_net_4;
wire   [3:0]     OE_DATA_81_const_net_4;
wire   [3:0]     OE_DATA_82_const_net_4;
wire   [3:0]     OE_DATA_83_const_net_4;
wire   [3:0]     OE_DATA_84_const_net_4;
wire   [3:0]     OE_DATA_85_const_net_4;
wire   [3:0]     OE_DATA_86_const_net_4;
wire   [3:0]     OE_DATA_87_const_net_4;
wire   [3:0]     OE_DATA_88_const_net_4;
wire   [3:0]     OE_DATA_89_const_net_4;
wire   [3:0]     OE_DATA_90_const_net_4;
wire   [3:0]     OE_DATA_91_const_net_4;
wire   [3:0]     OE_DATA_92_const_net_4;
wire   [3:0]     OE_DATA_93_const_net_4;
wire   [3:0]     OE_DATA_94_const_net_4;
wire   [3:0]     OE_DATA_95_const_net_4;
wire   [3:0]     OE_DATA_96_const_net_4;
wire   [3:0]     OE_DATA_97_const_net_4;
wire   [3:0]     OE_DATA_98_const_net_4;
wire   [3:0]     OE_DATA_99_const_net_4;
wire   [3:0]     OE_DATA_100_const_net_4;
wire   [3:0]     OE_DATA_101_const_net_4;
wire   [3:0]     OE_DATA_102_const_net_4;
wire   [3:0]     OE_DATA_103_const_net_4;
wire   [3:0]     OE_DATA_104_const_net_4;
wire   [3:0]     OE_DATA_105_const_net_4;
wire   [3:0]     OE_DATA_106_const_net_4;
wire   [3:0]     OE_DATA_107_const_net_4;
wire   [3:0]     OE_DATA_108_const_net_4;
wire   [3:0]     OE_DATA_109_const_net_4;
wire   [3:0]     OE_DATA_110_const_net_4;
wire   [3:0]     OE_DATA_111_const_net_4;
wire   [3:0]     OE_DATA_112_const_net_4;
wire   [3:0]     OE_DATA_113_const_net_4;
wire   [3:0]     OE_DATA_114_const_net_4;
wire   [3:0]     OE_DATA_115_const_net_4;
wire   [3:0]     OE_DATA_116_const_net_4;
wire   [3:0]     OE_DATA_117_const_net_4;
wire   [3:0]     OE_DATA_118_const_net_4;
wire   [3:0]     OE_DATA_119_const_net_4;
wire   [3:0]     OE_DATA_120_const_net_4;
wire   [3:0]     OE_DATA_121_const_net_4;
wire   [3:0]     OE_DATA_122_const_net_4;
wire   [3:0]     OE_DATA_123_const_net_4;
wire   [3:0]     OE_DATA_124_const_net_4;
wire   [3:0]     OE_DATA_125_const_net_4;
wire   [3:0]     OE_DATA_126_const_net_4;
wire   [3:0]     OE_DATA_127_const_net_4;
wire   [1:0]     PAD_const_net_1;
wire   [1:0]     PAD_I_const_net_1;
wire   [1:0]     PAD_N_const_net_1;
wire   [1:0]     PAD_I_N_const_net_1;
wire   [1:0]     RX_DQS_90_const_net_5;
wire   [2:0]     FIFO_WR_PTR_const_net_5;
wire   [2:0]     FIFO_RD_PTR_const_net_5;
wire   [2:0]     EYE_MONITOR_LANE_WIDTH_const_net_5;
wire   [7:0]     TX_DATA_0_const_net_8;
wire   [7:0]     TX_DATA_1_const_net_3;
wire   [7:0]     TX_DATA_2_const_net_4;
wire   [7:0]     TX_DATA_3_const_net_4;
wire   [7:0]     TX_DATA_4_const_net_4;
wire   [7:0]     TX_DATA_5_const_net_4;
wire   [7:0]     TX_DATA_6_const_net_4;
wire   [7:0]     TX_DATA_7_const_net_4;
wire   [7:0]     TX_DATA_8_const_net_4;
wire   [7:0]     TX_DATA_9_const_net_4;
wire   [7:0]     TX_DATA_10_const_net_4;
wire   [7:0]     TX_DATA_11_const_net_4;
wire   [7:0]     TX_DATA_12_const_net_5;
wire   [7:0]     TX_DATA_13_const_net_5;
wire   [7:0]     TX_DATA_14_const_net_5;
wire   [7:0]     TX_DATA_15_const_net_5;
wire   [7:0]     TX_DATA_16_const_net_5;
wire   [7:0]     TX_DATA_17_const_net_5;
wire   [7:0]     TX_DATA_18_const_net_5;
wire   [7:0]     TX_DATA_19_const_net_5;
wire   [7:0]     TX_DATA_20_const_net_5;
wire   [7:0]     TX_DATA_21_const_net_5;
wire   [7:0]     TX_DATA_22_const_net_5;
wire   [7:0]     TX_DATA_23_const_net_5;
wire   [7:0]     TX_DATA_24_const_net_5;
wire   [7:0]     TX_DATA_25_const_net_5;
wire   [7:0]     TX_DATA_26_const_net_5;
wire   [7:0]     TX_DATA_27_const_net_5;
wire   [7:0]     TX_DATA_28_const_net_5;
wire   [7:0]     TX_DATA_29_const_net_5;
wire   [7:0]     TX_DATA_30_const_net_5;
wire   [7:0]     TX_DATA_31_const_net_5;
wire   [7:0]     TX_DATA_32_const_net_5;
wire   [7:0]     TX_DATA_33_const_net_5;
wire   [7:0]     TX_DATA_34_const_net_5;
wire   [7:0]     TX_DATA_35_const_net_5;
wire   [7:0]     TX_DATA_36_const_net_5;
wire   [7:0]     TX_DATA_37_const_net_5;
wire   [7:0]     TX_DATA_38_const_net_5;
wire   [7:0]     TX_DATA_39_const_net_5;
wire   [7:0]     TX_DATA_40_const_net_5;
wire   [7:0]     TX_DATA_41_const_net_5;
wire   [7:0]     TX_DATA_42_const_net_5;
wire   [7:0]     TX_DATA_43_const_net_5;
wire   [7:0]     TX_DATA_44_const_net_5;
wire   [7:0]     TX_DATA_45_const_net_5;
wire   [7:0]     TX_DATA_46_const_net_5;
wire   [7:0]     TX_DATA_47_const_net_5;
wire   [7:0]     TX_DATA_48_const_net_5;
wire   [7:0]     TX_DATA_49_const_net_5;
wire   [7:0]     TX_DATA_50_const_net_5;
wire   [7:0]     TX_DATA_51_const_net_5;
wire   [7:0]     TX_DATA_52_const_net_5;
wire   [7:0]     TX_DATA_53_const_net_5;
wire   [7:0]     TX_DATA_54_const_net_5;
wire   [7:0]     TX_DATA_55_const_net_5;
wire   [7:0]     TX_DATA_56_const_net_5;
wire   [7:0]     TX_DATA_57_const_net_5;
wire   [7:0]     TX_DATA_58_const_net_5;
wire   [7:0]     TX_DATA_59_const_net_5;
wire   [7:0]     TX_DATA_60_const_net_5;
wire   [7:0]     TX_DATA_61_const_net_5;
wire   [7:0]     TX_DATA_62_const_net_5;
wire   [7:0]     TX_DATA_63_const_net_5;
wire   [7:0]     TX_DATA_64_const_net_5;
wire   [7:0]     TX_DATA_65_const_net_5;
wire   [7:0]     TX_DATA_66_const_net_5;
wire   [7:0]     TX_DATA_67_const_net_5;
wire   [7:0]     TX_DATA_68_const_net_5;
wire   [7:0]     TX_DATA_69_const_net_5;
wire   [7:0]     TX_DATA_70_const_net_5;
wire   [7:0]     TX_DATA_71_const_net_5;
wire   [7:0]     TX_DATA_72_const_net_5;
wire   [7:0]     TX_DATA_73_const_net_5;
wire   [7:0]     TX_DATA_74_const_net_5;
wire   [7:0]     TX_DATA_75_const_net_5;
wire   [7:0]     TX_DATA_76_const_net_5;
wire   [7:0]     TX_DATA_77_const_net_5;
wire   [7:0]     TX_DATA_78_const_net_5;
wire   [7:0]     TX_DATA_79_const_net_5;
wire   [7:0]     TX_DATA_80_const_net_5;
wire   [7:0]     TX_DATA_81_const_net_5;
wire   [7:0]     TX_DATA_82_const_net_5;
wire   [7:0]     TX_DATA_83_const_net_5;
wire   [7:0]     TX_DATA_84_const_net_5;
wire   [7:0]     TX_DATA_85_const_net_5;
wire   [7:0]     TX_DATA_86_const_net_5;
wire   [7:0]     TX_DATA_87_const_net_5;
wire   [7:0]     TX_DATA_88_const_net_5;
wire   [7:0]     TX_DATA_89_const_net_5;
wire   [7:0]     TX_DATA_90_const_net_5;
wire   [7:0]     TX_DATA_91_const_net_5;
wire   [7:0]     TX_DATA_92_const_net_5;
wire   [7:0]     TX_DATA_93_const_net_5;
wire   [7:0]     TX_DATA_94_const_net_5;
wire   [7:0]     TX_DATA_95_const_net_5;
wire   [7:0]     TX_DATA_96_const_net_5;
wire   [7:0]     TX_DATA_97_const_net_5;
wire   [7:0]     TX_DATA_98_const_net_5;
wire   [7:0]     TX_DATA_99_const_net_5;
wire   [7:0]     TX_DATA_100_const_net_5;
wire   [7:0]     TX_DATA_101_const_net_5;
wire   [7:0]     TX_DATA_102_const_net_5;
wire   [7:0]     TX_DATA_103_const_net_5;
wire   [7:0]     TX_DATA_104_const_net_5;
wire   [7:0]     TX_DATA_105_const_net_5;
wire   [7:0]     TX_DATA_106_const_net_5;
wire   [7:0]     TX_DATA_107_const_net_5;
wire   [7:0]     TX_DATA_108_const_net_5;
wire   [7:0]     TX_DATA_109_const_net_5;
wire   [7:0]     TX_DATA_110_const_net_5;
wire   [7:0]     TX_DATA_111_const_net_5;
wire   [7:0]     TX_DATA_112_const_net_5;
wire   [7:0]     TX_DATA_113_const_net_5;
wire   [7:0]     TX_DATA_114_const_net_5;
wire   [7:0]     TX_DATA_115_const_net_5;
wire   [7:0]     TX_DATA_116_const_net_5;
wire   [7:0]     TX_DATA_117_const_net_5;
wire   [7:0]     TX_DATA_118_const_net_5;
wire   [7:0]     TX_DATA_119_const_net_5;
wire   [7:0]     TX_DATA_120_const_net_5;
wire   [7:0]     TX_DATA_121_const_net_5;
wire   [7:0]     TX_DATA_122_const_net_5;
wire   [7:0]     TX_DATA_123_const_net_5;
wire   [7:0]     TX_DATA_124_const_net_5;
wire   [7:0]     TX_DATA_125_const_net_5;
wire   [7:0]     TX_DATA_126_const_net_5;
wire   [7:0]     TX_DATA_127_const_net_5;
wire   [3:0]     OE_DATA_0_const_net_16;
wire   [3:0]     OE_DATA_1_const_net_6;
wire   [3:0]     OE_DATA_2_const_net_5;
wire   [3:0]     OE_DATA_3_const_net_5;
wire   [3:0]     OE_DATA_4_const_net_5;
wire   [3:0]     OE_DATA_5_const_net_5;
wire   [3:0]     OE_DATA_6_const_net_5;
wire   [3:0]     OE_DATA_7_const_net_5;
wire   [3:0]     OE_DATA_8_const_net_5;
wire   [3:0]     OE_DATA_9_const_net_5;
wire   [3:0]     OE_DATA_10_const_net_5;
wire   [3:0]     OE_DATA_11_const_net_5;
wire   [3:0]     OE_DATA_12_const_net_5;
wire   [3:0]     OE_DATA_13_const_net_5;
wire   [3:0]     OE_DATA_14_const_net_5;
wire   [3:0]     OE_DATA_15_const_net_5;
wire   [3:0]     OE_DATA_16_const_net_5;
wire   [3:0]     OE_DATA_17_const_net_5;
wire   [3:0]     OE_DATA_18_const_net_5;
wire   [3:0]     OE_DATA_19_const_net_5;
wire   [3:0]     OE_DATA_20_const_net_5;
wire   [3:0]     OE_DATA_21_const_net_5;
wire   [3:0]     OE_DATA_22_const_net_5;
wire   [3:0]     OE_DATA_23_const_net_5;
wire   [3:0]     OE_DATA_24_const_net_5;
wire   [3:0]     OE_DATA_25_const_net_5;
wire   [3:0]     OE_DATA_26_const_net_5;
wire   [3:0]     OE_DATA_27_const_net_5;
wire   [3:0]     OE_DATA_28_const_net_5;
wire   [3:0]     OE_DATA_29_const_net_5;
wire   [3:0]     OE_DATA_30_const_net_5;
wire   [3:0]     OE_DATA_31_const_net_5;
wire   [3:0]     OE_DATA_32_const_net_5;
wire   [3:0]     OE_DATA_33_const_net_5;
wire   [3:0]     OE_DATA_34_const_net_5;
wire   [3:0]     OE_DATA_35_const_net_5;
wire   [3:0]     OE_DATA_36_const_net_5;
wire   [3:0]     OE_DATA_37_const_net_5;
wire   [3:0]     OE_DATA_38_const_net_5;
wire   [3:0]     OE_DATA_39_const_net_5;
wire   [3:0]     OE_DATA_40_const_net_5;
wire   [3:0]     OE_DATA_41_const_net_5;
wire   [3:0]     OE_DATA_42_const_net_5;
wire   [3:0]     OE_DATA_43_const_net_5;
wire   [3:0]     OE_DATA_44_const_net_5;
wire   [3:0]     OE_DATA_45_const_net_5;
wire   [3:0]     OE_DATA_46_const_net_5;
wire   [3:0]     OE_DATA_47_const_net_5;
wire   [3:0]     OE_DATA_48_const_net_5;
wire   [3:0]     OE_DATA_49_const_net_5;
wire   [3:0]     OE_DATA_50_const_net_5;
wire   [3:0]     OE_DATA_51_const_net_5;
wire   [3:0]     OE_DATA_52_const_net_5;
wire   [3:0]     OE_DATA_53_const_net_5;
wire   [3:0]     OE_DATA_54_const_net_5;
wire   [3:0]     OE_DATA_55_const_net_5;
wire   [3:0]     OE_DATA_56_const_net_5;
wire   [3:0]     OE_DATA_57_const_net_5;
wire   [3:0]     OE_DATA_58_const_net_5;
wire   [3:0]     OE_DATA_59_const_net_5;
wire   [3:0]     OE_DATA_60_const_net_5;
wire   [3:0]     OE_DATA_61_const_net_5;
wire   [3:0]     OE_DATA_62_const_net_5;
wire   [3:0]     OE_DATA_63_const_net_5;
wire   [3:0]     OE_DATA_64_const_net_5;
wire   [3:0]     OE_DATA_65_const_net_5;
wire   [3:0]     OE_DATA_66_const_net_5;
wire   [3:0]     OE_DATA_67_const_net_5;
wire   [3:0]     OE_DATA_68_const_net_5;
wire   [3:0]     OE_DATA_69_const_net_5;
wire   [3:0]     OE_DATA_70_const_net_5;
wire   [3:0]     OE_DATA_71_const_net_5;
wire   [3:0]     OE_DATA_72_const_net_5;
wire   [3:0]     OE_DATA_73_const_net_5;
wire   [3:0]     OE_DATA_74_const_net_5;
wire   [3:0]     OE_DATA_75_const_net_5;
wire   [3:0]     OE_DATA_76_const_net_5;
wire   [3:0]     OE_DATA_77_const_net_5;
wire   [3:0]     OE_DATA_78_const_net_5;
wire   [3:0]     OE_DATA_79_const_net_5;
wire   [3:0]     OE_DATA_80_const_net_5;
wire   [3:0]     OE_DATA_81_const_net_5;
wire   [3:0]     OE_DATA_82_const_net_5;
wire   [3:0]     OE_DATA_83_const_net_5;
wire   [3:0]     OE_DATA_84_const_net_5;
wire   [3:0]     OE_DATA_85_const_net_5;
wire   [3:0]     OE_DATA_86_const_net_5;
wire   [3:0]     OE_DATA_87_const_net_5;
wire   [3:0]     OE_DATA_88_const_net_5;
wire   [3:0]     OE_DATA_89_const_net_5;
wire   [3:0]     OE_DATA_90_const_net_5;
wire   [3:0]     OE_DATA_91_const_net_5;
wire   [3:0]     OE_DATA_92_const_net_5;
wire   [3:0]     OE_DATA_93_const_net_5;
wire   [3:0]     OE_DATA_94_const_net_5;
wire   [3:0]     OE_DATA_95_const_net_5;
wire   [3:0]     OE_DATA_96_const_net_5;
wire   [3:0]     OE_DATA_97_const_net_5;
wire   [3:0]     OE_DATA_98_const_net_5;
wire   [3:0]     OE_DATA_99_const_net_5;
wire   [3:0]     OE_DATA_100_const_net_5;
wire   [3:0]     OE_DATA_101_const_net_5;
wire   [3:0]     OE_DATA_102_const_net_5;
wire   [3:0]     OE_DATA_103_const_net_5;
wire   [3:0]     OE_DATA_104_const_net_5;
wire   [3:0]     OE_DATA_105_const_net_5;
wire   [3:0]     OE_DATA_106_const_net_5;
wire   [3:0]     OE_DATA_107_const_net_5;
wire   [3:0]     OE_DATA_108_const_net_5;
wire   [3:0]     OE_DATA_109_const_net_5;
wire   [3:0]     OE_DATA_110_const_net_5;
wire   [3:0]     OE_DATA_111_const_net_5;
wire   [3:0]     OE_DATA_112_const_net_5;
wire   [3:0]     OE_DATA_113_const_net_5;
wire   [3:0]     OE_DATA_114_const_net_5;
wire   [3:0]     OE_DATA_115_const_net_5;
wire   [3:0]     OE_DATA_116_const_net_5;
wire   [3:0]     OE_DATA_117_const_net_5;
wire   [3:0]     OE_DATA_118_const_net_5;
wire   [3:0]     OE_DATA_119_const_net_5;
wire   [3:0]     OE_DATA_120_const_net_5;
wire   [3:0]     OE_DATA_121_const_net_5;
wire   [3:0]     OE_DATA_122_const_net_5;
wire   [3:0]     OE_DATA_123_const_net_5;
wire   [3:0]     OE_DATA_124_const_net_5;
wire   [3:0]     OE_DATA_125_const_net_5;
wire   [3:0]     OE_DATA_126_const_net_5;
wire   [3:0]     OE_DATA_127_const_net_5;
wire   [1:0]     RX_DQS_90_const_net_6;
wire   [2:0]     FIFO_WR_PTR_const_net_6;
wire   [2:0]     FIFO_RD_PTR_const_net_6;
wire   [2:0]     EYE_MONITOR_LANE_WIDTH_const_net_6;
wire   [3:0]     TX_DATA_2_const_net_5;
wire   [3:0]     TX_DATA_3_const_net_5;
wire   [3:0]     TX_DATA_4_const_net_5;
wire   [3:0]     TX_DATA_5_const_net_5;
wire   [3:0]     TX_DATA_6_const_net_5;
wire   [3:0]     TX_DATA_7_const_net_5;
wire   [3:0]     TX_DATA_8_const_net_5;
wire   [3:0]     TX_DATA_9_const_net_5;
wire   [3:0]     TX_DATA_10_const_net_5;
wire   [3:0]     TX_DATA_11_const_net_5;
wire   [3:0]     TX_DATA_12_const_net_6;
wire   [3:0]     TX_DATA_13_const_net_6;
wire   [3:0]     TX_DATA_14_const_net_6;
wire   [3:0]     TX_DATA_15_const_net_6;
wire   [3:0]     TX_DATA_16_const_net_6;
wire   [3:0]     TX_DATA_17_const_net_6;
wire   [3:0]     TX_DATA_18_const_net_6;
wire   [3:0]     TX_DATA_19_const_net_6;
wire   [3:0]     TX_DATA_20_const_net_6;
wire   [3:0]     TX_DATA_21_const_net_6;
wire   [3:0]     TX_DATA_22_const_net_6;
wire   [3:0]     TX_DATA_23_const_net_6;
wire   [3:0]     TX_DATA_24_const_net_6;
wire   [3:0]     TX_DATA_25_const_net_6;
wire   [3:0]     TX_DATA_26_const_net_6;
wire   [3:0]     TX_DATA_27_const_net_6;
wire   [3:0]     TX_DATA_28_const_net_6;
wire   [3:0]     TX_DATA_29_const_net_6;
wire   [3:0]     TX_DATA_30_const_net_6;
wire   [3:0]     TX_DATA_31_const_net_6;
wire   [3:0]     TX_DATA_32_const_net_6;
wire   [3:0]     TX_DATA_33_const_net_6;
wire   [3:0]     TX_DATA_34_const_net_6;
wire   [3:0]     TX_DATA_35_const_net_6;
wire   [3:0]     TX_DATA_36_const_net_6;
wire   [3:0]     TX_DATA_37_const_net_6;
wire   [3:0]     TX_DATA_38_const_net_6;
wire   [3:0]     TX_DATA_39_const_net_6;
wire   [3:0]     TX_DATA_40_const_net_6;
wire   [3:0]     TX_DATA_41_const_net_6;
wire   [3:0]     TX_DATA_42_const_net_6;
wire   [3:0]     TX_DATA_43_const_net_6;
wire   [3:0]     TX_DATA_44_const_net_6;
wire   [3:0]     TX_DATA_45_const_net_6;
wire   [3:0]     TX_DATA_46_const_net_6;
wire   [3:0]     TX_DATA_47_const_net_6;
wire   [3:0]     TX_DATA_48_const_net_6;
wire   [3:0]     TX_DATA_49_const_net_6;
wire   [3:0]     TX_DATA_50_const_net_6;
wire   [3:0]     TX_DATA_51_const_net_6;
wire   [3:0]     TX_DATA_52_const_net_6;
wire   [3:0]     TX_DATA_53_const_net_6;
wire   [3:0]     TX_DATA_54_const_net_6;
wire   [3:0]     TX_DATA_55_const_net_6;
wire   [3:0]     TX_DATA_56_const_net_6;
wire   [3:0]     TX_DATA_57_const_net_6;
wire   [3:0]     TX_DATA_58_const_net_6;
wire   [3:0]     TX_DATA_59_const_net_6;
wire   [3:0]     TX_DATA_60_const_net_6;
wire   [3:0]     TX_DATA_61_const_net_6;
wire   [3:0]     TX_DATA_62_const_net_6;
wire   [3:0]     TX_DATA_63_const_net_6;
wire   [3:0]     TX_DATA_64_const_net_6;
wire   [3:0]     TX_DATA_65_const_net_6;
wire   [3:0]     TX_DATA_66_const_net_6;
wire   [3:0]     TX_DATA_67_const_net_6;
wire   [3:0]     TX_DATA_68_const_net_6;
wire   [3:0]     TX_DATA_69_const_net_6;
wire   [3:0]     TX_DATA_70_const_net_6;
wire   [3:0]     TX_DATA_71_const_net_6;
wire   [3:0]     TX_DATA_72_const_net_6;
wire   [3:0]     TX_DATA_73_const_net_6;
wire   [3:0]     TX_DATA_74_const_net_6;
wire   [3:0]     TX_DATA_75_const_net_6;
wire   [3:0]     TX_DATA_76_const_net_6;
wire   [3:0]     TX_DATA_77_const_net_6;
wire   [3:0]     TX_DATA_78_const_net_6;
wire   [3:0]     TX_DATA_79_const_net_6;
wire   [3:0]     TX_DATA_80_const_net_6;
wire   [3:0]     TX_DATA_81_const_net_6;
wire   [3:0]     TX_DATA_82_const_net_6;
wire   [3:0]     TX_DATA_83_const_net_6;
wire   [3:0]     TX_DATA_84_const_net_6;
wire   [3:0]     TX_DATA_85_const_net_6;
wire   [3:0]     TX_DATA_86_const_net_6;
wire   [3:0]     TX_DATA_87_const_net_6;
wire   [3:0]     TX_DATA_88_const_net_6;
wire   [3:0]     TX_DATA_89_const_net_6;
wire   [3:0]     TX_DATA_90_const_net_6;
wire   [3:0]     TX_DATA_91_const_net_6;
wire   [3:0]     TX_DATA_92_const_net_6;
wire   [3:0]     TX_DATA_93_const_net_6;
wire   [3:0]     TX_DATA_94_const_net_6;
wire   [3:0]     TX_DATA_95_const_net_6;
wire   [3:0]     TX_DATA_96_const_net_6;
wire   [3:0]     TX_DATA_97_const_net_6;
wire   [3:0]     TX_DATA_98_const_net_6;
wire   [3:0]     TX_DATA_99_const_net_6;
wire   [3:0]     TX_DATA_100_const_net_6;
wire   [3:0]     TX_DATA_101_const_net_6;
wire   [3:0]     TX_DATA_102_const_net_6;
wire   [3:0]     TX_DATA_103_const_net_6;
wire   [3:0]     TX_DATA_104_const_net_6;
wire   [3:0]     TX_DATA_105_const_net_6;
wire   [3:0]     TX_DATA_106_const_net_6;
wire   [3:0]     TX_DATA_107_const_net_6;
wire   [3:0]     TX_DATA_108_const_net_6;
wire   [3:0]     TX_DATA_109_const_net_6;
wire   [3:0]     TX_DATA_110_const_net_6;
wire   [3:0]     TX_DATA_111_const_net_6;
wire   [3:0]     TX_DATA_112_const_net_6;
wire   [3:0]     TX_DATA_113_const_net_6;
wire   [3:0]     TX_DATA_114_const_net_6;
wire   [3:0]     TX_DATA_115_const_net_6;
wire   [3:0]     TX_DATA_116_const_net_6;
wire   [3:0]     TX_DATA_117_const_net_6;
wire   [3:0]     TX_DATA_118_const_net_6;
wire   [3:0]     TX_DATA_119_const_net_6;
wire   [3:0]     TX_DATA_120_const_net_6;
wire   [3:0]     TX_DATA_121_const_net_6;
wire   [3:0]     TX_DATA_122_const_net_6;
wire   [3:0]     TX_DATA_123_const_net_6;
wire   [3:0]     TX_DATA_124_const_net_6;
wire   [3:0]     TX_DATA_125_const_net_6;
wire   [3:0]     TX_DATA_126_const_net_6;
wire   [3:0]     TX_DATA_127_const_net_6;
wire   [3:0]     OE_DATA_2_const_net_6;
wire   [3:0]     OE_DATA_3_const_net_6;
wire   [3:0]     OE_DATA_4_const_net_6;
wire   [3:0]     OE_DATA_5_const_net_6;
wire   [3:0]     OE_DATA_6_const_net_6;
wire   [3:0]     OE_DATA_7_const_net_6;
wire   [3:0]     OE_DATA_8_const_net_6;
wire   [3:0]     OE_DATA_9_const_net_6;
wire   [3:0]     OE_DATA_10_const_net_6;
wire   [3:0]     OE_DATA_11_const_net_6;
wire   [3:0]     OE_DATA_12_const_net_6;
wire   [3:0]     OE_DATA_13_const_net_6;
wire   [3:0]     OE_DATA_14_const_net_6;
wire   [3:0]     OE_DATA_15_const_net_6;
wire   [3:0]     OE_DATA_16_const_net_6;
wire   [3:0]     OE_DATA_17_const_net_6;
wire   [3:0]     OE_DATA_18_const_net_6;
wire   [3:0]     OE_DATA_19_const_net_6;
wire   [3:0]     OE_DATA_20_const_net_6;
wire   [3:0]     OE_DATA_21_const_net_6;
wire   [3:0]     OE_DATA_22_const_net_6;
wire   [3:0]     OE_DATA_23_const_net_6;
wire   [3:0]     OE_DATA_24_const_net_6;
wire   [3:0]     OE_DATA_25_const_net_6;
wire   [3:0]     OE_DATA_26_const_net_6;
wire   [3:0]     OE_DATA_27_const_net_6;
wire   [3:0]     OE_DATA_28_const_net_6;
wire   [3:0]     OE_DATA_29_const_net_6;
wire   [3:0]     OE_DATA_30_const_net_6;
wire   [3:0]     OE_DATA_31_const_net_6;
wire   [3:0]     OE_DATA_32_const_net_6;
wire   [3:0]     OE_DATA_33_const_net_6;
wire   [3:0]     OE_DATA_34_const_net_6;
wire   [3:0]     OE_DATA_35_const_net_6;
wire   [3:0]     OE_DATA_36_const_net_6;
wire   [3:0]     OE_DATA_37_const_net_6;
wire   [3:0]     OE_DATA_38_const_net_6;
wire   [3:0]     OE_DATA_39_const_net_6;
wire   [3:0]     OE_DATA_40_const_net_6;
wire   [3:0]     OE_DATA_41_const_net_6;
wire   [3:0]     OE_DATA_42_const_net_6;
wire   [3:0]     OE_DATA_43_const_net_6;
wire   [3:0]     OE_DATA_44_const_net_6;
wire   [3:0]     OE_DATA_45_const_net_6;
wire   [3:0]     OE_DATA_46_const_net_6;
wire   [3:0]     OE_DATA_47_const_net_6;
wire   [3:0]     OE_DATA_48_const_net_6;
wire   [3:0]     OE_DATA_49_const_net_6;
wire   [3:0]     OE_DATA_50_const_net_6;
wire   [3:0]     OE_DATA_51_const_net_6;
wire   [3:0]     OE_DATA_52_const_net_6;
wire   [3:0]     OE_DATA_53_const_net_6;
wire   [3:0]     OE_DATA_54_const_net_6;
wire   [3:0]     OE_DATA_55_const_net_6;
wire   [3:0]     OE_DATA_56_const_net_6;
wire   [3:0]     OE_DATA_57_const_net_6;
wire   [3:0]     OE_DATA_58_const_net_6;
wire   [3:0]     OE_DATA_59_const_net_6;
wire   [3:0]     OE_DATA_60_const_net_6;
wire   [3:0]     OE_DATA_61_const_net_6;
wire   [3:0]     OE_DATA_62_const_net_6;
wire   [3:0]     OE_DATA_63_const_net_6;
wire   [3:0]     OE_DATA_64_const_net_6;
wire   [3:0]     OE_DATA_65_const_net_6;
wire   [3:0]     OE_DATA_66_const_net_6;
wire   [3:0]     OE_DATA_67_const_net_6;
wire   [3:0]     OE_DATA_68_const_net_6;
wire   [3:0]     OE_DATA_69_const_net_6;
wire   [3:0]     OE_DATA_70_const_net_6;
wire   [3:0]     OE_DATA_71_const_net_6;
wire   [3:0]     OE_DATA_72_const_net_6;
wire   [3:0]     OE_DATA_73_const_net_6;
wire   [3:0]     OE_DATA_74_const_net_6;
wire   [3:0]     OE_DATA_75_const_net_6;
wire   [3:0]     OE_DATA_76_const_net_6;
wire   [3:0]     OE_DATA_77_const_net_6;
wire   [3:0]     OE_DATA_78_const_net_6;
wire   [3:0]     OE_DATA_79_const_net_6;
wire   [3:0]     OE_DATA_80_const_net_6;
wire   [3:0]     OE_DATA_81_const_net_6;
wire   [3:0]     OE_DATA_82_const_net_6;
wire   [3:0]     OE_DATA_83_const_net_6;
wire   [3:0]     OE_DATA_84_const_net_6;
wire   [3:0]     OE_DATA_85_const_net_6;
wire   [3:0]     OE_DATA_86_const_net_6;
wire   [3:0]     OE_DATA_87_const_net_6;
wire   [3:0]     OE_DATA_88_const_net_6;
wire   [3:0]     OE_DATA_89_const_net_6;
wire   [3:0]     OE_DATA_90_const_net_6;
wire   [3:0]     OE_DATA_91_const_net_6;
wire   [3:0]     OE_DATA_92_const_net_6;
wire   [3:0]     OE_DATA_93_const_net_6;
wire   [3:0]     OE_DATA_94_const_net_6;
wire   [3:0]     OE_DATA_95_const_net_6;
wire   [3:0]     OE_DATA_96_const_net_6;
wire   [3:0]     OE_DATA_97_const_net_6;
wire   [3:0]     OE_DATA_98_const_net_6;
wire   [3:0]     OE_DATA_99_const_net_6;
wire   [3:0]     OE_DATA_100_const_net_6;
wire   [3:0]     OE_DATA_101_const_net_6;
wire   [3:0]     OE_DATA_102_const_net_6;
wire   [3:0]     OE_DATA_103_const_net_6;
wire   [3:0]     OE_DATA_104_const_net_6;
wire   [3:0]     OE_DATA_105_const_net_6;
wire   [3:0]     OE_DATA_106_const_net_6;
wire   [3:0]     OE_DATA_107_const_net_6;
wire   [3:0]     OE_DATA_108_const_net_6;
wire   [3:0]     OE_DATA_109_const_net_6;
wire   [3:0]     OE_DATA_110_const_net_6;
wire   [3:0]     OE_DATA_111_const_net_6;
wire   [3:0]     OE_DATA_112_const_net_6;
wire   [3:0]     OE_DATA_113_const_net_6;
wire   [3:0]     OE_DATA_114_const_net_6;
wire   [3:0]     OE_DATA_115_const_net_6;
wire   [3:0]     OE_DATA_116_const_net_6;
wire   [3:0]     OE_DATA_117_const_net_6;
wire   [3:0]     OE_DATA_118_const_net_6;
wire   [3:0]     OE_DATA_119_const_net_6;
wire   [3:0]     OE_DATA_120_const_net_6;
wire   [3:0]     OE_DATA_121_const_net_6;
wire   [3:0]     OE_DATA_122_const_net_6;
wire   [3:0]     OE_DATA_123_const_net_6;
wire   [3:0]     OE_DATA_124_const_net_6;
wire   [3:0]     OE_DATA_125_const_net_6;
wire   [3:0]     OE_DATA_126_const_net_6;
wire   [3:0]     OE_DATA_127_const_net_6;
wire   [1:0]     PAD_const_net_2;
wire   [1:0]     PAD_I_const_net_2;
wire   [1:0]     PAD_N_const_net_2;
wire   [1:0]     PAD_I_N_const_net_2;
wire   [1:0]     RX_DQS_90_const_net_7;
wire   [2:0]     FIFO_WR_PTR_const_net_7;
wire   [2:0]     FIFO_RD_PTR_const_net_7;
wire   [2:0]     EYE_MONITOR_LANE_WIDTH_const_net_7;
wire   [3:0]     TX_DATA_1_const_net_4;
wire   [3:0]     TX_DATA_2_const_net_6;
wire   [3:0]     TX_DATA_3_const_net_6;
wire   [3:0]     TX_DATA_4_const_net_6;
wire   [3:0]     TX_DATA_5_const_net_6;
wire   [3:0]     TX_DATA_6_const_net_6;
wire   [3:0]     TX_DATA_7_const_net_6;
wire   [3:0]     TX_DATA_8_const_net_6;
wire   [3:0]     TX_DATA_9_const_net_6;
wire   [3:0]     TX_DATA_10_const_net_6;
wire   [3:0]     TX_DATA_11_const_net_6;
wire   [3:0]     TX_DATA_12_const_net_7;
wire   [3:0]     TX_DATA_13_const_net_7;
wire   [3:0]     TX_DATA_14_const_net_7;
wire   [3:0]     TX_DATA_15_const_net_7;
wire   [3:0]     TX_DATA_16_const_net_7;
wire   [3:0]     TX_DATA_17_const_net_7;
wire   [3:0]     TX_DATA_18_const_net_7;
wire   [3:0]     TX_DATA_19_const_net_7;
wire   [3:0]     TX_DATA_20_const_net_7;
wire   [3:0]     TX_DATA_21_const_net_7;
wire   [3:0]     TX_DATA_22_const_net_7;
wire   [3:0]     TX_DATA_23_const_net_7;
wire   [3:0]     TX_DATA_24_const_net_7;
wire   [3:0]     TX_DATA_25_const_net_7;
wire   [3:0]     TX_DATA_26_const_net_7;
wire   [3:0]     TX_DATA_27_const_net_7;
wire   [3:0]     TX_DATA_28_const_net_7;
wire   [3:0]     TX_DATA_29_const_net_7;
wire   [3:0]     TX_DATA_30_const_net_7;
wire   [3:0]     TX_DATA_31_const_net_7;
wire   [3:0]     TX_DATA_32_const_net_7;
wire   [3:0]     TX_DATA_33_const_net_7;
wire   [3:0]     TX_DATA_34_const_net_7;
wire   [3:0]     TX_DATA_35_const_net_7;
wire   [3:0]     TX_DATA_36_const_net_7;
wire   [3:0]     TX_DATA_37_const_net_7;
wire   [3:0]     TX_DATA_38_const_net_7;
wire   [3:0]     TX_DATA_39_const_net_7;
wire   [3:0]     TX_DATA_40_const_net_7;
wire   [3:0]     TX_DATA_41_const_net_7;
wire   [3:0]     TX_DATA_42_const_net_7;
wire   [3:0]     TX_DATA_43_const_net_7;
wire   [3:0]     TX_DATA_44_const_net_7;
wire   [3:0]     TX_DATA_45_const_net_7;
wire   [3:0]     TX_DATA_46_const_net_7;
wire   [3:0]     TX_DATA_47_const_net_7;
wire   [3:0]     TX_DATA_48_const_net_7;
wire   [3:0]     TX_DATA_49_const_net_7;
wire   [3:0]     TX_DATA_50_const_net_7;
wire   [3:0]     TX_DATA_51_const_net_7;
wire   [3:0]     TX_DATA_52_const_net_7;
wire   [3:0]     TX_DATA_53_const_net_7;
wire   [3:0]     TX_DATA_54_const_net_7;
wire   [3:0]     TX_DATA_55_const_net_7;
wire   [3:0]     TX_DATA_56_const_net_7;
wire   [3:0]     TX_DATA_57_const_net_7;
wire   [3:0]     TX_DATA_58_const_net_7;
wire   [3:0]     TX_DATA_59_const_net_7;
wire   [3:0]     TX_DATA_60_const_net_7;
wire   [3:0]     TX_DATA_61_const_net_7;
wire   [3:0]     TX_DATA_62_const_net_7;
wire   [3:0]     TX_DATA_63_const_net_7;
wire   [3:0]     TX_DATA_64_const_net_7;
wire   [3:0]     TX_DATA_65_const_net_7;
wire   [3:0]     TX_DATA_66_const_net_7;
wire   [3:0]     TX_DATA_67_const_net_7;
wire   [3:0]     TX_DATA_68_const_net_7;
wire   [3:0]     TX_DATA_69_const_net_7;
wire   [3:0]     TX_DATA_70_const_net_7;
wire   [3:0]     TX_DATA_71_const_net_7;
wire   [3:0]     TX_DATA_72_const_net_7;
wire   [3:0]     TX_DATA_73_const_net_7;
wire   [3:0]     TX_DATA_74_const_net_7;
wire   [3:0]     TX_DATA_75_const_net_7;
wire   [3:0]     TX_DATA_76_const_net_7;
wire   [3:0]     TX_DATA_77_const_net_7;
wire   [3:0]     TX_DATA_78_const_net_7;
wire   [3:0]     TX_DATA_79_const_net_7;
wire   [3:0]     TX_DATA_80_const_net_7;
wire   [3:0]     TX_DATA_81_const_net_7;
wire   [3:0]     TX_DATA_82_const_net_7;
wire   [3:0]     TX_DATA_83_const_net_7;
wire   [3:0]     TX_DATA_84_const_net_7;
wire   [3:0]     TX_DATA_85_const_net_7;
wire   [3:0]     TX_DATA_86_const_net_7;
wire   [3:0]     TX_DATA_87_const_net_7;
wire   [3:0]     TX_DATA_88_const_net_7;
wire   [3:0]     TX_DATA_89_const_net_7;
wire   [3:0]     TX_DATA_90_const_net_7;
wire   [3:0]     TX_DATA_91_const_net_7;
wire   [3:0]     TX_DATA_92_const_net_7;
wire   [3:0]     TX_DATA_93_const_net_7;
wire   [3:0]     TX_DATA_94_const_net_7;
wire   [3:0]     TX_DATA_95_const_net_7;
wire   [3:0]     TX_DATA_96_const_net_7;
wire   [3:0]     TX_DATA_97_const_net_7;
wire   [3:0]     TX_DATA_98_const_net_7;
wire   [3:0]     TX_DATA_99_const_net_7;
wire   [3:0]     TX_DATA_100_const_net_7;
wire   [3:0]     TX_DATA_101_const_net_7;
wire   [3:0]     TX_DATA_102_const_net_7;
wire   [3:0]     TX_DATA_103_const_net_7;
wire   [3:0]     TX_DATA_104_const_net_7;
wire   [3:0]     TX_DATA_105_const_net_7;
wire   [3:0]     TX_DATA_106_const_net_7;
wire   [3:0]     TX_DATA_107_const_net_7;
wire   [3:0]     TX_DATA_108_const_net_7;
wire   [3:0]     TX_DATA_109_const_net_7;
wire   [3:0]     TX_DATA_110_const_net_7;
wire   [3:0]     TX_DATA_111_const_net_7;
wire   [3:0]     TX_DATA_112_const_net_7;
wire   [3:0]     TX_DATA_113_const_net_7;
wire   [3:0]     TX_DATA_114_const_net_7;
wire   [3:0]     TX_DATA_115_const_net_7;
wire   [3:0]     TX_DATA_116_const_net_7;
wire   [3:0]     TX_DATA_117_const_net_7;
wire   [3:0]     TX_DATA_118_const_net_7;
wire   [3:0]     TX_DATA_119_const_net_7;
wire   [3:0]     TX_DATA_120_const_net_7;
wire   [3:0]     TX_DATA_121_const_net_7;
wire   [3:0]     TX_DATA_122_const_net_7;
wire   [3:0]     TX_DATA_123_const_net_7;
wire   [3:0]     TX_DATA_124_const_net_7;
wire   [3:0]     TX_DATA_125_const_net_7;
wire   [3:0]     TX_DATA_126_const_net_7;
wire   [3:0]     TX_DATA_127_const_net_7;
wire   [3:0]     OE_DATA_1_const_net_7;
wire   [3:0]     OE_DATA_2_const_net_7;
wire   [3:0]     OE_DATA_3_const_net_7;
wire   [3:0]     OE_DATA_4_const_net_7;
wire   [3:0]     OE_DATA_5_const_net_7;
wire   [3:0]     OE_DATA_6_const_net_7;
wire   [3:0]     OE_DATA_7_const_net_7;
wire   [3:0]     OE_DATA_8_const_net_7;
wire   [3:0]     OE_DATA_9_const_net_7;
wire   [3:0]     OE_DATA_10_const_net_7;
wire   [3:0]     OE_DATA_11_const_net_7;
wire   [3:0]     OE_DATA_12_const_net_7;
wire   [3:0]     OE_DATA_13_const_net_7;
wire   [3:0]     OE_DATA_14_const_net_7;
wire   [3:0]     OE_DATA_15_const_net_7;
wire   [3:0]     OE_DATA_16_const_net_7;
wire   [3:0]     OE_DATA_17_const_net_7;
wire   [3:0]     OE_DATA_18_const_net_7;
wire   [3:0]     OE_DATA_19_const_net_7;
wire   [3:0]     OE_DATA_20_const_net_7;
wire   [3:0]     OE_DATA_21_const_net_7;
wire   [3:0]     OE_DATA_22_const_net_7;
wire   [3:0]     OE_DATA_23_const_net_7;
wire   [3:0]     OE_DATA_24_const_net_7;
wire   [3:0]     OE_DATA_25_const_net_7;
wire   [3:0]     OE_DATA_26_const_net_7;
wire   [3:0]     OE_DATA_27_const_net_7;
wire   [3:0]     OE_DATA_28_const_net_7;
wire   [3:0]     OE_DATA_29_const_net_7;
wire   [3:0]     OE_DATA_30_const_net_7;
wire   [3:0]     OE_DATA_31_const_net_7;
wire   [3:0]     OE_DATA_32_const_net_7;
wire   [3:0]     OE_DATA_33_const_net_7;
wire   [3:0]     OE_DATA_34_const_net_7;
wire   [3:0]     OE_DATA_35_const_net_7;
wire   [3:0]     OE_DATA_36_const_net_7;
wire   [3:0]     OE_DATA_37_const_net_7;
wire   [3:0]     OE_DATA_38_const_net_7;
wire   [3:0]     OE_DATA_39_const_net_7;
wire   [3:0]     OE_DATA_40_const_net_7;
wire   [3:0]     OE_DATA_41_const_net_7;
wire   [3:0]     OE_DATA_42_const_net_7;
wire   [3:0]     OE_DATA_43_const_net_7;
wire   [3:0]     OE_DATA_44_const_net_7;
wire   [3:0]     OE_DATA_45_const_net_7;
wire   [3:0]     OE_DATA_46_const_net_7;
wire   [3:0]     OE_DATA_47_const_net_7;
wire   [3:0]     OE_DATA_48_const_net_7;
wire   [3:0]     OE_DATA_49_const_net_7;
wire   [3:0]     OE_DATA_50_const_net_7;
wire   [3:0]     OE_DATA_51_const_net_7;
wire   [3:0]     OE_DATA_52_const_net_7;
wire   [3:0]     OE_DATA_53_const_net_7;
wire   [3:0]     OE_DATA_54_const_net_7;
wire   [3:0]     OE_DATA_55_const_net_7;
wire   [3:0]     OE_DATA_56_const_net_7;
wire   [3:0]     OE_DATA_57_const_net_7;
wire   [3:0]     OE_DATA_58_const_net_7;
wire   [3:0]     OE_DATA_59_const_net_7;
wire   [3:0]     OE_DATA_60_const_net_7;
wire   [3:0]     OE_DATA_61_const_net_7;
wire   [3:0]     OE_DATA_62_const_net_7;
wire   [3:0]     OE_DATA_63_const_net_7;
wire   [3:0]     OE_DATA_64_const_net_7;
wire   [3:0]     OE_DATA_65_const_net_7;
wire   [3:0]     OE_DATA_66_const_net_7;
wire   [3:0]     OE_DATA_67_const_net_7;
wire   [3:0]     OE_DATA_68_const_net_7;
wire   [3:0]     OE_DATA_69_const_net_7;
wire   [3:0]     OE_DATA_70_const_net_7;
wire   [3:0]     OE_DATA_71_const_net_7;
wire   [3:0]     OE_DATA_72_const_net_7;
wire   [3:0]     OE_DATA_73_const_net_7;
wire   [3:0]     OE_DATA_74_const_net_7;
wire   [3:0]     OE_DATA_75_const_net_7;
wire   [3:0]     OE_DATA_76_const_net_7;
wire   [3:0]     OE_DATA_77_const_net_7;
wire   [3:0]     OE_DATA_78_const_net_7;
wire   [3:0]     OE_DATA_79_const_net_7;
wire   [3:0]     OE_DATA_80_const_net_7;
wire   [3:0]     OE_DATA_81_const_net_7;
wire   [3:0]     OE_DATA_82_const_net_7;
wire   [3:0]     OE_DATA_83_const_net_7;
wire   [3:0]     OE_DATA_84_const_net_7;
wire   [3:0]     OE_DATA_85_const_net_7;
wire   [3:0]     OE_DATA_86_const_net_7;
wire   [3:0]     OE_DATA_87_const_net_7;
wire   [3:0]     OE_DATA_88_const_net_7;
wire   [3:0]     OE_DATA_89_const_net_7;
wire   [3:0]     OE_DATA_90_const_net_7;
wire   [3:0]     OE_DATA_91_const_net_7;
wire   [3:0]     OE_DATA_92_const_net_7;
wire   [3:0]     OE_DATA_93_const_net_7;
wire   [3:0]     OE_DATA_94_const_net_7;
wire   [3:0]     OE_DATA_95_const_net_7;
wire   [3:0]     OE_DATA_96_const_net_7;
wire   [3:0]     OE_DATA_97_const_net_7;
wire   [3:0]     OE_DATA_98_const_net_7;
wire   [3:0]     OE_DATA_99_const_net_7;
wire   [3:0]     OE_DATA_100_const_net_7;
wire   [3:0]     OE_DATA_101_const_net_7;
wire   [3:0]     OE_DATA_102_const_net_7;
wire   [3:0]     OE_DATA_103_const_net_7;
wire   [3:0]     OE_DATA_104_const_net_7;
wire   [3:0]     OE_DATA_105_const_net_7;
wire   [3:0]     OE_DATA_106_const_net_7;
wire   [3:0]     OE_DATA_107_const_net_7;
wire   [3:0]     OE_DATA_108_const_net_7;
wire   [3:0]     OE_DATA_109_const_net_7;
wire   [3:0]     OE_DATA_110_const_net_7;
wire   [3:0]     OE_DATA_111_const_net_7;
wire   [3:0]     OE_DATA_112_const_net_7;
wire   [3:0]     OE_DATA_113_const_net_7;
wire   [3:0]     OE_DATA_114_const_net_7;
wire   [3:0]     OE_DATA_115_const_net_7;
wire   [3:0]     OE_DATA_116_const_net_7;
wire   [3:0]     OE_DATA_117_const_net_7;
wire   [3:0]     OE_DATA_118_const_net_7;
wire   [3:0]     OE_DATA_119_const_net_7;
wire   [3:0]     OE_DATA_120_const_net_7;
wire   [3:0]     OE_DATA_121_const_net_7;
wire   [3:0]     OE_DATA_122_const_net_7;
wire   [3:0]     OE_DATA_123_const_net_7;
wire   [3:0]     OE_DATA_124_const_net_7;
wire   [3:0]     OE_DATA_125_const_net_7;
wire   [3:0]     OE_DATA_126_const_net_7;
wire   [3:0]     OE_DATA_127_const_net_7;
wire   [1:0]     RX_DQS_90_const_net_8;
wire   [2:0]     FIFO_WR_PTR_const_net_8;
wire   [2:0]     FIFO_RD_PTR_const_net_8;
wire   [2:0]     EYE_MONITOR_LANE_WIDTH_const_net_8;
wire   [3:0]     TX_DATA_1_const_net_5;
wire   [3:0]     TX_DATA_2_const_net_7;
wire   [3:0]     TX_DATA_3_const_net_7;
wire   [3:0]     TX_DATA_4_const_net_7;
wire   [3:0]     TX_DATA_5_const_net_7;
wire   [3:0]     TX_DATA_6_const_net_7;
wire   [3:0]     TX_DATA_7_const_net_7;
wire   [3:0]     TX_DATA_8_const_net_7;
wire   [3:0]     TX_DATA_9_const_net_7;
wire   [3:0]     TX_DATA_10_const_net_7;
wire   [3:0]     TX_DATA_11_const_net_7;
wire   [3:0]     TX_DATA_12_const_net_8;
wire   [3:0]     TX_DATA_13_const_net_8;
wire   [3:0]     TX_DATA_14_const_net_8;
wire   [3:0]     TX_DATA_15_const_net_8;
wire   [3:0]     TX_DATA_16_const_net_8;
wire   [3:0]     TX_DATA_17_const_net_8;
wire   [3:0]     TX_DATA_18_const_net_8;
wire   [3:0]     TX_DATA_19_const_net_8;
wire   [3:0]     TX_DATA_20_const_net_8;
wire   [3:0]     TX_DATA_21_const_net_8;
wire   [3:0]     TX_DATA_22_const_net_8;
wire   [3:0]     TX_DATA_23_const_net_8;
wire   [3:0]     TX_DATA_24_const_net_8;
wire   [3:0]     TX_DATA_25_const_net_8;
wire   [3:0]     TX_DATA_26_const_net_8;
wire   [3:0]     TX_DATA_27_const_net_8;
wire   [3:0]     TX_DATA_28_const_net_8;
wire   [3:0]     TX_DATA_29_const_net_8;
wire   [3:0]     TX_DATA_30_const_net_8;
wire   [3:0]     TX_DATA_31_const_net_8;
wire   [3:0]     TX_DATA_32_const_net_8;
wire   [3:0]     TX_DATA_33_const_net_8;
wire   [3:0]     TX_DATA_34_const_net_8;
wire   [3:0]     TX_DATA_35_const_net_8;
wire   [3:0]     TX_DATA_36_const_net_8;
wire   [3:0]     TX_DATA_37_const_net_8;
wire   [3:0]     TX_DATA_38_const_net_8;
wire   [3:0]     TX_DATA_39_const_net_8;
wire   [3:0]     TX_DATA_40_const_net_8;
wire   [3:0]     TX_DATA_41_const_net_8;
wire   [3:0]     TX_DATA_42_const_net_8;
wire   [3:0]     TX_DATA_43_const_net_8;
wire   [3:0]     TX_DATA_44_const_net_8;
wire   [3:0]     TX_DATA_45_const_net_8;
wire   [3:0]     TX_DATA_46_const_net_8;
wire   [3:0]     TX_DATA_47_const_net_8;
wire   [3:0]     TX_DATA_48_const_net_8;
wire   [3:0]     TX_DATA_49_const_net_8;
wire   [3:0]     TX_DATA_50_const_net_8;
wire   [3:0]     TX_DATA_51_const_net_8;
wire   [3:0]     TX_DATA_52_const_net_8;
wire   [3:0]     TX_DATA_53_const_net_8;
wire   [3:0]     TX_DATA_54_const_net_8;
wire   [3:0]     TX_DATA_55_const_net_8;
wire   [3:0]     TX_DATA_56_const_net_8;
wire   [3:0]     TX_DATA_57_const_net_8;
wire   [3:0]     TX_DATA_58_const_net_8;
wire   [3:0]     TX_DATA_59_const_net_8;
wire   [3:0]     TX_DATA_60_const_net_8;
wire   [3:0]     TX_DATA_61_const_net_8;
wire   [3:0]     TX_DATA_62_const_net_8;
wire   [3:0]     TX_DATA_63_const_net_8;
wire   [3:0]     TX_DATA_64_const_net_8;
wire   [3:0]     TX_DATA_65_const_net_8;
wire   [3:0]     TX_DATA_66_const_net_8;
wire   [3:0]     TX_DATA_67_const_net_8;
wire   [3:0]     TX_DATA_68_const_net_8;
wire   [3:0]     TX_DATA_69_const_net_8;
wire   [3:0]     TX_DATA_70_const_net_8;
wire   [3:0]     TX_DATA_71_const_net_8;
wire   [3:0]     TX_DATA_72_const_net_8;
wire   [3:0]     TX_DATA_73_const_net_8;
wire   [3:0]     TX_DATA_74_const_net_8;
wire   [3:0]     TX_DATA_75_const_net_8;
wire   [3:0]     TX_DATA_76_const_net_8;
wire   [3:0]     TX_DATA_77_const_net_8;
wire   [3:0]     TX_DATA_78_const_net_8;
wire   [3:0]     TX_DATA_79_const_net_8;
wire   [3:0]     TX_DATA_80_const_net_8;
wire   [3:0]     TX_DATA_81_const_net_8;
wire   [3:0]     TX_DATA_82_const_net_8;
wire   [3:0]     TX_DATA_83_const_net_8;
wire   [3:0]     TX_DATA_84_const_net_8;
wire   [3:0]     TX_DATA_85_const_net_8;
wire   [3:0]     TX_DATA_86_const_net_8;
wire   [3:0]     TX_DATA_87_const_net_8;
wire   [3:0]     TX_DATA_88_const_net_8;
wire   [3:0]     TX_DATA_89_const_net_8;
wire   [3:0]     TX_DATA_90_const_net_8;
wire   [3:0]     TX_DATA_91_const_net_8;
wire   [3:0]     TX_DATA_92_const_net_8;
wire   [3:0]     TX_DATA_93_const_net_8;
wire   [3:0]     TX_DATA_94_const_net_8;
wire   [3:0]     TX_DATA_95_const_net_8;
wire   [3:0]     TX_DATA_96_const_net_8;
wire   [3:0]     TX_DATA_97_const_net_8;
wire   [3:0]     TX_DATA_98_const_net_8;
wire   [3:0]     TX_DATA_99_const_net_8;
wire   [3:0]     TX_DATA_100_const_net_8;
wire   [3:0]     TX_DATA_101_const_net_8;
wire   [3:0]     TX_DATA_102_const_net_8;
wire   [3:0]     TX_DATA_103_const_net_8;
wire   [3:0]     TX_DATA_104_const_net_8;
wire   [3:0]     TX_DATA_105_const_net_8;
wire   [3:0]     TX_DATA_106_const_net_8;
wire   [3:0]     TX_DATA_107_const_net_8;
wire   [3:0]     TX_DATA_108_const_net_8;
wire   [3:0]     TX_DATA_109_const_net_8;
wire   [3:0]     TX_DATA_110_const_net_8;
wire   [3:0]     TX_DATA_111_const_net_8;
wire   [3:0]     TX_DATA_112_const_net_8;
wire   [3:0]     TX_DATA_113_const_net_8;
wire   [3:0]     TX_DATA_114_const_net_8;
wire   [3:0]     TX_DATA_115_const_net_8;
wire   [3:0]     TX_DATA_116_const_net_8;
wire   [3:0]     TX_DATA_117_const_net_8;
wire   [3:0]     TX_DATA_118_const_net_8;
wire   [3:0]     TX_DATA_119_const_net_8;
wire   [3:0]     TX_DATA_120_const_net_8;
wire   [3:0]     TX_DATA_121_const_net_8;
wire   [3:0]     TX_DATA_122_const_net_8;
wire   [3:0]     TX_DATA_123_const_net_8;
wire   [3:0]     TX_DATA_124_const_net_8;
wire   [3:0]     TX_DATA_125_const_net_8;
wire   [3:0]     TX_DATA_126_const_net_8;
wire   [3:0]     TX_DATA_127_const_net_8;
wire   [3:0]     OE_DATA_1_const_net_8;
wire   [3:0]     OE_DATA_2_const_net_8;
wire   [3:0]     OE_DATA_3_const_net_8;
wire   [3:0]     OE_DATA_4_const_net_8;
wire   [3:0]     OE_DATA_5_const_net_8;
wire   [3:0]     OE_DATA_6_const_net_8;
wire   [3:0]     OE_DATA_7_const_net_8;
wire   [3:0]     OE_DATA_8_const_net_8;
wire   [3:0]     OE_DATA_9_const_net_8;
wire   [3:0]     OE_DATA_10_const_net_8;
wire   [3:0]     OE_DATA_11_const_net_8;
wire   [3:0]     OE_DATA_12_const_net_8;
wire   [3:0]     OE_DATA_13_const_net_8;
wire   [3:0]     OE_DATA_14_const_net_8;
wire   [3:0]     OE_DATA_15_const_net_8;
wire   [3:0]     OE_DATA_16_const_net_8;
wire   [3:0]     OE_DATA_17_const_net_8;
wire   [3:0]     OE_DATA_18_const_net_8;
wire   [3:0]     OE_DATA_19_const_net_8;
wire   [3:0]     OE_DATA_20_const_net_8;
wire   [3:0]     OE_DATA_21_const_net_8;
wire   [3:0]     OE_DATA_22_const_net_8;
wire   [3:0]     OE_DATA_23_const_net_8;
wire   [3:0]     OE_DATA_24_const_net_8;
wire   [3:0]     OE_DATA_25_const_net_8;
wire   [3:0]     OE_DATA_26_const_net_8;
wire   [3:0]     OE_DATA_27_const_net_8;
wire   [3:0]     OE_DATA_28_const_net_8;
wire   [3:0]     OE_DATA_29_const_net_8;
wire   [3:0]     OE_DATA_30_const_net_8;
wire   [3:0]     OE_DATA_31_const_net_8;
wire   [3:0]     OE_DATA_32_const_net_8;
wire   [3:0]     OE_DATA_33_const_net_8;
wire   [3:0]     OE_DATA_34_const_net_8;
wire   [3:0]     OE_DATA_35_const_net_8;
wire   [3:0]     OE_DATA_36_const_net_8;
wire   [3:0]     OE_DATA_37_const_net_8;
wire   [3:0]     OE_DATA_38_const_net_8;
wire   [3:0]     OE_DATA_39_const_net_8;
wire   [3:0]     OE_DATA_40_const_net_8;
wire   [3:0]     OE_DATA_41_const_net_8;
wire   [3:0]     OE_DATA_42_const_net_8;
wire   [3:0]     OE_DATA_43_const_net_8;
wire   [3:0]     OE_DATA_44_const_net_8;
wire   [3:0]     OE_DATA_45_const_net_8;
wire   [3:0]     OE_DATA_46_const_net_8;
wire   [3:0]     OE_DATA_47_const_net_8;
wire   [3:0]     OE_DATA_48_const_net_8;
wire   [3:0]     OE_DATA_49_const_net_8;
wire   [3:0]     OE_DATA_50_const_net_8;
wire   [3:0]     OE_DATA_51_const_net_8;
wire   [3:0]     OE_DATA_52_const_net_8;
wire   [3:0]     OE_DATA_53_const_net_8;
wire   [3:0]     OE_DATA_54_const_net_8;
wire   [3:0]     OE_DATA_55_const_net_8;
wire   [3:0]     OE_DATA_56_const_net_8;
wire   [3:0]     OE_DATA_57_const_net_8;
wire   [3:0]     OE_DATA_58_const_net_8;
wire   [3:0]     OE_DATA_59_const_net_8;
wire   [3:0]     OE_DATA_60_const_net_8;
wire   [3:0]     OE_DATA_61_const_net_8;
wire   [3:0]     OE_DATA_62_const_net_8;
wire   [3:0]     OE_DATA_63_const_net_8;
wire   [3:0]     OE_DATA_64_const_net_8;
wire   [3:0]     OE_DATA_65_const_net_8;
wire   [3:0]     OE_DATA_66_const_net_8;
wire   [3:0]     OE_DATA_67_const_net_8;
wire   [3:0]     OE_DATA_68_const_net_8;
wire   [3:0]     OE_DATA_69_const_net_8;
wire   [3:0]     OE_DATA_70_const_net_8;
wire   [3:0]     OE_DATA_71_const_net_8;
wire   [3:0]     OE_DATA_72_const_net_8;
wire   [3:0]     OE_DATA_73_const_net_8;
wire   [3:0]     OE_DATA_74_const_net_8;
wire   [3:0]     OE_DATA_75_const_net_8;
wire   [3:0]     OE_DATA_76_const_net_8;
wire   [3:0]     OE_DATA_77_const_net_8;
wire   [3:0]     OE_DATA_78_const_net_8;
wire   [3:0]     OE_DATA_79_const_net_8;
wire   [3:0]     OE_DATA_80_const_net_8;
wire   [3:0]     OE_DATA_81_const_net_8;
wire   [3:0]     OE_DATA_82_const_net_8;
wire   [3:0]     OE_DATA_83_const_net_8;
wire   [3:0]     OE_DATA_84_const_net_8;
wire   [3:0]     OE_DATA_85_const_net_8;
wire   [3:0]     OE_DATA_86_const_net_8;
wire   [3:0]     OE_DATA_87_const_net_8;
wire   [3:0]     OE_DATA_88_const_net_8;
wire   [3:0]     OE_DATA_89_const_net_8;
wire   [3:0]     OE_DATA_90_const_net_8;
wire   [3:0]     OE_DATA_91_const_net_8;
wire   [3:0]     OE_DATA_92_const_net_8;
wire   [3:0]     OE_DATA_93_const_net_8;
wire   [3:0]     OE_DATA_94_const_net_8;
wire   [3:0]     OE_DATA_95_const_net_8;
wire   [3:0]     OE_DATA_96_const_net_8;
wire   [3:0]     OE_DATA_97_const_net_8;
wire   [3:0]     OE_DATA_98_const_net_8;
wire   [3:0]     OE_DATA_99_const_net_8;
wire   [3:0]     OE_DATA_100_const_net_8;
wire   [3:0]     OE_DATA_101_const_net_8;
wire   [3:0]     OE_DATA_102_const_net_8;
wire   [3:0]     OE_DATA_103_const_net_8;
wire   [3:0]     OE_DATA_104_const_net_8;
wire   [3:0]     OE_DATA_105_const_net_8;
wire   [3:0]     OE_DATA_106_const_net_8;
wire   [3:0]     OE_DATA_107_const_net_8;
wire   [3:0]     OE_DATA_108_const_net_8;
wire   [3:0]     OE_DATA_109_const_net_8;
wire   [3:0]     OE_DATA_110_const_net_8;
wire   [3:0]     OE_DATA_111_const_net_8;
wire   [3:0]     OE_DATA_112_const_net_8;
wire   [3:0]     OE_DATA_113_const_net_8;
wire   [3:0]     OE_DATA_114_const_net_8;
wire   [3:0]     OE_DATA_115_const_net_8;
wire   [3:0]     OE_DATA_116_const_net_8;
wire   [3:0]     OE_DATA_117_const_net_8;
wire   [3:0]     OE_DATA_118_const_net_8;
wire   [3:0]     OE_DATA_119_const_net_8;
wire   [3:0]     OE_DATA_120_const_net_8;
wire   [3:0]     OE_DATA_121_const_net_8;
wire   [3:0]     OE_DATA_122_const_net_8;
wire   [3:0]     OE_DATA_123_const_net_8;
wire   [3:0]     OE_DATA_124_const_net_8;
wire   [3:0]     OE_DATA_125_const_net_8;
wire   [3:0]     OE_DATA_126_const_net_8;
wire   [3:0]     OE_DATA_127_const_net_8;
wire   [1:0]     RX_DQS_90_const_net_9;
wire   [2:0]     FIFO_WR_PTR_const_net_9;
wire   [2:0]     FIFO_RD_PTR_const_net_9;
wire   [2:0]     EYE_MONITOR_LANE_WIDTH_const_net_9;
wire   [3:0]     TX_DATA_1_const_net_6;
wire   [3:0]     TX_DATA_2_const_net_8;
wire   [3:0]     TX_DATA_3_const_net_8;
wire   [3:0]     TX_DATA_4_const_net_8;
wire   [3:0]     TX_DATA_5_const_net_8;
wire   [3:0]     TX_DATA_6_const_net_8;
wire   [3:0]     TX_DATA_7_const_net_8;
wire   [3:0]     TX_DATA_8_const_net_8;
wire   [3:0]     TX_DATA_9_const_net_8;
wire   [3:0]     TX_DATA_10_const_net_8;
wire   [3:0]     TX_DATA_11_const_net_8;
wire   [3:0]     TX_DATA_12_const_net_9;
wire   [3:0]     TX_DATA_13_const_net_9;
wire   [3:0]     TX_DATA_14_const_net_9;
wire   [3:0]     TX_DATA_15_const_net_9;
wire   [3:0]     TX_DATA_16_const_net_9;
wire   [3:0]     TX_DATA_17_const_net_9;
wire   [3:0]     TX_DATA_18_const_net_9;
wire   [3:0]     TX_DATA_19_const_net_9;
wire   [3:0]     TX_DATA_20_const_net_9;
wire   [3:0]     TX_DATA_21_const_net_9;
wire   [3:0]     TX_DATA_22_const_net_9;
wire   [3:0]     TX_DATA_23_const_net_9;
wire   [3:0]     TX_DATA_24_const_net_9;
wire   [3:0]     TX_DATA_25_const_net_9;
wire   [3:0]     TX_DATA_26_const_net_9;
wire   [3:0]     TX_DATA_27_const_net_9;
wire   [3:0]     TX_DATA_28_const_net_9;
wire   [3:0]     TX_DATA_29_const_net_9;
wire   [3:0]     TX_DATA_30_const_net_9;
wire   [3:0]     TX_DATA_31_const_net_9;
wire   [3:0]     TX_DATA_32_const_net_9;
wire   [3:0]     TX_DATA_33_const_net_9;
wire   [3:0]     TX_DATA_34_const_net_9;
wire   [3:0]     TX_DATA_35_const_net_9;
wire   [3:0]     TX_DATA_36_const_net_9;
wire   [3:0]     TX_DATA_37_const_net_9;
wire   [3:0]     TX_DATA_38_const_net_9;
wire   [3:0]     TX_DATA_39_const_net_9;
wire   [3:0]     TX_DATA_40_const_net_9;
wire   [3:0]     TX_DATA_41_const_net_9;
wire   [3:0]     TX_DATA_42_const_net_9;
wire   [3:0]     TX_DATA_43_const_net_9;
wire   [3:0]     TX_DATA_44_const_net_9;
wire   [3:0]     TX_DATA_45_const_net_9;
wire   [3:0]     TX_DATA_46_const_net_9;
wire   [3:0]     TX_DATA_47_const_net_9;
wire   [3:0]     TX_DATA_48_const_net_9;
wire   [3:0]     TX_DATA_49_const_net_9;
wire   [3:0]     TX_DATA_50_const_net_9;
wire   [3:0]     TX_DATA_51_const_net_9;
wire   [3:0]     TX_DATA_52_const_net_9;
wire   [3:0]     TX_DATA_53_const_net_9;
wire   [3:0]     TX_DATA_54_const_net_9;
wire   [3:0]     TX_DATA_55_const_net_9;
wire   [3:0]     TX_DATA_56_const_net_9;
wire   [3:0]     TX_DATA_57_const_net_9;
wire   [3:0]     TX_DATA_58_const_net_9;
wire   [3:0]     TX_DATA_59_const_net_9;
wire   [3:0]     TX_DATA_60_const_net_9;
wire   [3:0]     TX_DATA_61_const_net_9;
wire   [3:0]     TX_DATA_62_const_net_9;
wire   [3:0]     TX_DATA_63_const_net_9;
wire   [3:0]     TX_DATA_64_const_net_9;
wire   [3:0]     TX_DATA_65_const_net_9;
wire   [3:0]     TX_DATA_66_const_net_9;
wire   [3:0]     TX_DATA_67_const_net_9;
wire   [3:0]     TX_DATA_68_const_net_9;
wire   [3:0]     TX_DATA_69_const_net_9;
wire   [3:0]     TX_DATA_70_const_net_9;
wire   [3:0]     TX_DATA_71_const_net_9;
wire   [3:0]     TX_DATA_72_const_net_9;
wire   [3:0]     TX_DATA_73_const_net_9;
wire   [3:0]     TX_DATA_74_const_net_9;
wire   [3:0]     TX_DATA_75_const_net_9;
wire   [3:0]     TX_DATA_76_const_net_9;
wire   [3:0]     TX_DATA_77_const_net_9;
wire   [3:0]     TX_DATA_78_const_net_9;
wire   [3:0]     TX_DATA_79_const_net_9;
wire   [3:0]     TX_DATA_80_const_net_9;
wire   [3:0]     TX_DATA_81_const_net_9;
wire   [3:0]     TX_DATA_82_const_net_9;
wire   [3:0]     TX_DATA_83_const_net_9;
wire   [3:0]     TX_DATA_84_const_net_9;
wire   [3:0]     TX_DATA_85_const_net_9;
wire   [3:0]     TX_DATA_86_const_net_9;
wire   [3:0]     TX_DATA_87_const_net_9;
wire   [3:0]     TX_DATA_88_const_net_9;
wire   [3:0]     TX_DATA_89_const_net_9;
wire   [3:0]     TX_DATA_90_const_net_9;
wire   [3:0]     TX_DATA_91_const_net_9;
wire   [3:0]     TX_DATA_92_const_net_9;
wire   [3:0]     TX_DATA_93_const_net_9;
wire   [3:0]     TX_DATA_94_const_net_9;
wire   [3:0]     TX_DATA_95_const_net_9;
wire   [3:0]     TX_DATA_96_const_net_9;
wire   [3:0]     TX_DATA_97_const_net_9;
wire   [3:0]     TX_DATA_98_const_net_9;
wire   [3:0]     TX_DATA_99_const_net_9;
wire   [3:0]     TX_DATA_100_const_net_9;
wire   [3:0]     TX_DATA_101_const_net_9;
wire   [3:0]     TX_DATA_102_const_net_9;
wire   [3:0]     TX_DATA_103_const_net_9;
wire   [3:0]     TX_DATA_104_const_net_9;
wire   [3:0]     TX_DATA_105_const_net_9;
wire   [3:0]     TX_DATA_106_const_net_9;
wire   [3:0]     TX_DATA_107_const_net_9;
wire   [3:0]     TX_DATA_108_const_net_9;
wire   [3:0]     TX_DATA_109_const_net_9;
wire   [3:0]     TX_DATA_110_const_net_9;
wire   [3:0]     TX_DATA_111_const_net_9;
wire   [3:0]     TX_DATA_112_const_net_9;
wire   [3:0]     TX_DATA_113_const_net_9;
wire   [3:0]     TX_DATA_114_const_net_9;
wire   [3:0]     TX_DATA_115_const_net_9;
wire   [3:0]     TX_DATA_116_const_net_9;
wire   [3:0]     TX_DATA_117_const_net_9;
wire   [3:0]     TX_DATA_118_const_net_9;
wire   [3:0]     TX_DATA_119_const_net_9;
wire   [3:0]     TX_DATA_120_const_net_9;
wire   [3:0]     TX_DATA_121_const_net_9;
wire   [3:0]     TX_DATA_122_const_net_9;
wire   [3:0]     TX_DATA_123_const_net_9;
wire   [3:0]     TX_DATA_124_const_net_9;
wire   [3:0]     TX_DATA_125_const_net_9;
wire   [3:0]     TX_DATA_126_const_net_9;
wire   [3:0]     TX_DATA_127_const_net_9;
wire   [3:0]     OE_DATA_1_const_net_9;
wire   [3:0]     OE_DATA_2_const_net_9;
wire   [3:0]     OE_DATA_3_const_net_9;
wire   [3:0]     OE_DATA_4_const_net_9;
wire   [3:0]     OE_DATA_5_const_net_9;
wire   [3:0]     OE_DATA_6_const_net_9;
wire   [3:0]     OE_DATA_7_const_net_9;
wire   [3:0]     OE_DATA_8_const_net_9;
wire   [3:0]     OE_DATA_9_const_net_9;
wire   [3:0]     OE_DATA_10_const_net_9;
wire   [3:0]     OE_DATA_11_const_net_9;
wire   [3:0]     OE_DATA_12_const_net_9;
wire   [3:0]     OE_DATA_13_const_net_9;
wire   [3:0]     OE_DATA_14_const_net_9;
wire   [3:0]     OE_DATA_15_const_net_9;
wire   [3:0]     OE_DATA_16_const_net_9;
wire   [3:0]     OE_DATA_17_const_net_9;
wire   [3:0]     OE_DATA_18_const_net_9;
wire   [3:0]     OE_DATA_19_const_net_9;
wire   [3:0]     OE_DATA_20_const_net_9;
wire   [3:0]     OE_DATA_21_const_net_9;
wire   [3:0]     OE_DATA_22_const_net_9;
wire   [3:0]     OE_DATA_23_const_net_9;
wire   [3:0]     OE_DATA_24_const_net_9;
wire   [3:0]     OE_DATA_25_const_net_9;
wire   [3:0]     OE_DATA_26_const_net_9;
wire   [3:0]     OE_DATA_27_const_net_9;
wire   [3:0]     OE_DATA_28_const_net_9;
wire   [3:0]     OE_DATA_29_const_net_9;
wire   [3:0]     OE_DATA_30_const_net_9;
wire   [3:0]     OE_DATA_31_const_net_9;
wire   [3:0]     OE_DATA_32_const_net_9;
wire   [3:0]     OE_DATA_33_const_net_9;
wire   [3:0]     OE_DATA_34_const_net_9;
wire   [3:0]     OE_DATA_35_const_net_9;
wire   [3:0]     OE_DATA_36_const_net_9;
wire   [3:0]     OE_DATA_37_const_net_9;
wire   [3:0]     OE_DATA_38_const_net_9;
wire   [3:0]     OE_DATA_39_const_net_9;
wire   [3:0]     OE_DATA_40_const_net_9;
wire   [3:0]     OE_DATA_41_const_net_9;
wire   [3:0]     OE_DATA_42_const_net_9;
wire   [3:0]     OE_DATA_43_const_net_9;
wire   [3:0]     OE_DATA_44_const_net_9;
wire   [3:0]     OE_DATA_45_const_net_9;
wire   [3:0]     OE_DATA_46_const_net_9;
wire   [3:0]     OE_DATA_47_const_net_9;
wire   [3:0]     OE_DATA_48_const_net_9;
wire   [3:0]     OE_DATA_49_const_net_9;
wire   [3:0]     OE_DATA_50_const_net_9;
wire   [3:0]     OE_DATA_51_const_net_9;
wire   [3:0]     OE_DATA_52_const_net_9;
wire   [3:0]     OE_DATA_53_const_net_9;
wire   [3:0]     OE_DATA_54_const_net_9;
wire   [3:0]     OE_DATA_55_const_net_9;
wire   [3:0]     OE_DATA_56_const_net_9;
wire   [3:0]     OE_DATA_57_const_net_9;
wire   [3:0]     OE_DATA_58_const_net_9;
wire   [3:0]     OE_DATA_59_const_net_9;
wire   [3:0]     OE_DATA_60_const_net_9;
wire   [3:0]     OE_DATA_61_const_net_9;
wire   [3:0]     OE_DATA_62_const_net_9;
wire   [3:0]     OE_DATA_63_const_net_9;
wire   [3:0]     OE_DATA_64_const_net_9;
wire   [3:0]     OE_DATA_65_const_net_9;
wire   [3:0]     OE_DATA_66_const_net_9;
wire   [3:0]     OE_DATA_67_const_net_9;
wire   [3:0]     OE_DATA_68_const_net_9;
wire   [3:0]     OE_DATA_69_const_net_9;
wire   [3:0]     OE_DATA_70_const_net_9;
wire   [3:0]     OE_DATA_71_const_net_9;
wire   [3:0]     OE_DATA_72_const_net_9;
wire   [3:0]     OE_DATA_73_const_net_9;
wire   [3:0]     OE_DATA_74_const_net_9;
wire   [3:0]     OE_DATA_75_const_net_9;
wire   [3:0]     OE_DATA_76_const_net_9;
wire   [3:0]     OE_DATA_77_const_net_9;
wire   [3:0]     OE_DATA_78_const_net_9;
wire   [3:0]     OE_DATA_79_const_net_9;
wire   [3:0]     OE_DATA_80_const_net_9;
wire   [3:0]     OE_DATA_81_const_net_9;
wire   [3:0]     OE_DATA_82_const_net_9;
wire   [3:0]     OE_DATA_83_const_net_9;
wire   [3:0]     OE_DATA_84_const_net_9;
wire   [3:0]     OE_DATA_85_const_net_9;
wire   [3:0]     OE_DATA_86_const_net_9;
wire   [3:0]     OE_DATA_87_const_net_9;
wire   [3:0]     OE_DATA_88_const_net_9;
wire   [3:0]     OE_DATA_89_const_net_9;
wire   [3:0]     OE_DATA_90_const_net_9;
wire   [3:0]     OE_DATA_91_const_net_9;
wire   [3:0]     OE_DATA_92_const_net_9;
wire   [3:0]     OE_DATA_93_const_net_9;
wire   [3:0]     OE_DATA_94_const_net_9;
wire   [3:0]     OE_DATA_95_const_net_9;
wire   [3:0]     OE_DATA_96_const_net_9;
wire   [3:0]     OE_DATA_97_const_net_9;
wire   [3:0]     OE_DATA_98_const_net_9;
wire   [3:0]     OE_DATA_99_const_net_9;
wire   [3:0]     OE_DATA_100_const_net_9;
wire   [3:0]     OE_DATA_101_const_net_9;
wire   [3:0]     OE_DATA_102_const_net_9;
wire   [3:0]     OE_DATA_103_const_net_9;
wire   [3:0]     OE_DATA_104_const_net_9;
wire   [3:0]     OE_DATA_105_const_net_9;
wire   [3:0]     OE_DATA_106_const_net_9;
wire   [3:0]     OE_DATA_107_const_net_9;
wire   [3:0]     OE_DATA_108_const_net_9;
wire   [3:0]     OE_DATA_109_const_net_9;
wire   [3:0]     OE_DATA_110_const_net_9;
wire   [3:0]     OE_DATA_111_const_net_9;
wire   [3:0]     OE_DATA_112_const_net_9;
wire   [3:0]     OE_DATA_113_const_net_9;
wire   [3:0]     OE_DATA_114_const_net_9;
wire   [3:0]     OE_DATA_115_const_net_9;
wire   [3:0]     OE_DATA_116_const_net_9;
wire   [3:0]     OE_DATA_117_const_net_9;
wire   [3:0]     OE_DATA_118_const_net_9;
wire   [3:0]     OE_DATA_119_const_net_9;
wire   [3:0]     OE_DATA_120_const_net_9;
wire   [3:0]     OE_DATA_121_const_net_9;
wire   [3:0]     OE_DATA_122_const_net_9;
wire   [3:0]     OE_DATA_123_const_net_9;
wire   [3:0]     OE_DATA_124_const_net_9;
wire   [3:0]     OE_DATA_125_const_net_9;
wire   [3:0]     OE_DATA_126_const_net_9;
wire   [3:0]     OE_DATA_127_const_net_9;
wire   [1:0]     RX_DQS_90_const_net_10;
wire   [2:0]     FIFO_WR_PTR_const_net_10;
wire   [2:0]     FIFO_RD_PTR_const_net_10;
wire   [2:0]     EYE_MONITOR_LANE_WIDTH_const_net_10;
wire   [3:0]     TX_DATA_1_const_net_7;
wire   [3:0]     TX_DATA_2_const_net_9;
wire   [3:0]     TX_DATA_3_const_net_9;
wire   [3:0]     TX_DATA_4_const_net_9;
wire   [3:0]     TX_DATA_5_const_net_9;
wire   [3:0]     TX_DATA_6_const_net_9;
wire   [3:0]     TX_DATA_7_const_net_9;
wire   [3:0]     TX_DATA_8_const_net_9;
wire   [3:0]     TX_DATA_9_const_net_9;
wire   [3:0]     TX_DATA_10_const_net_9;
wire   [3:0]     TX_DATA_11_const_net_9;
wire   [3:0]     TX_DATA_12_const_net_10;
wire   [3:0]     TX_DATA_13_const_net_10;
wire   [3:0]     TX_DATA_14_const_net_10;
wire   [3:0]     TX_DATA_15_const_net_10;
wire   [3:0]     TX_DATA_16_const_net_10;
wire   [3:0]     TX_DATA_17_const_net_10;
wire   [3:0]     TX_DATA_18_const_net_10;
wire   [3:0]     TX_DATA_19_const_net_10;
wire   [3:0]     TX_DATA_20_const_net_10;
wire   [3:0]     TX_DATA_21_const_net_10;
wire   [3:0]     TX_DATA_22_const_net_10;
wire   [3:0]     TX_DATA_23_const_net_10;
wire   [3:0]     TX_DATA_24_const_net_10;
wire   [3:0]     TX_DATA_25_const_net_10;
wire   [3:0]     TX_DATA_26_const_net_10;
wire   [3:0]     TX_DATA_27_const_net_10;
wire   [3:0]     TX_DATA_28_const_net_10;
wire   [3:0]     TX_DATA_29_const_net_10;
wire   [3:0]     TX_DATA_30_const_net_10;
wire   [3:0]     TX_DATA_31_const_net_10;
wire   [3:0]     TX_DATA_32_const_net_10;
wire   [3:0]     TX_DATA_33_const_net_10;
wire   [3:0]     TX_DATA_34_const_net_10;
wire   [3:0]     TX_DATA_35_const_net_10;
wire   [3:0]     TX_DATA_36_const_net_10;
wire   [3:0]     TX_DATA_37_const_net_10;
wire   [3:0]     TX_DATA_38_const_net_10;
wire   [3:0]     TX_DATA_39_const_net_10;
wire   [3:0]     TX_DATA_40_const_net_10;
wire   [3:0]     TX_DATA_41_const_net_10;
wire   [3:0]     TX_DATA_42_const_net_10;
wire   [3:0]     TX_DATA_43_const_net_10;
wire   [3:0]     TX_DATA_44_const_net_10;
wire   [3:0]     TX_DATA_45_const_net_10;
wire   [3:0]     TX_DATA_46_const_net_10;
wire   [3:0]     TX_DATA_47_const_net_10;
wire   [3:0]     TX_DATA_48_const_net_10;
wire   [3:0]     TX_DATA_49_const_net_10;
wire   [3:0]     TX_DATA_50_const_net_10;
wire   [3:0]     TX_DATA_51_const_net_10;
wire   [3:0]     TX_DATA_52_const_net_10;
wire   [3:0]     TX_DATA_53_const_net_10;
wire   [3:0]     TX_DATA_54_const_net_10;
wire   [3:0]     TX_DATA_55_const_net_10;
wire   [3:0]     TX_DATA_56_const_net_10;
wire   [3:0]     TX_DATA_57_const_net_10;
wire   [3:0]     TX_DATA_58_const_net_10;
wire   [3:0]     TX_DATA_59_const_net_10;
wire   [3:0]     TX_DATA_60_const_net_10;
wire   [3:0]     TX_DATA_61_const_net_10;
wire   [3:0]     TX_DATA_62_const_net_10;
wire   [3:0]     TX_DATA_63_const_net_10;
wire   [3:0]     TX_DATA_64_const_net_10;
wire   [3:0]     TX_DATA_65_const_net_10;
wire   [3:0]     TX_DATA_66_const_net_10;
wire   [3:0]     TX_DATA_67_const_net_10;
wire   [3:0]     TX_DATA_68_const_net_10;
wire   [3:0]     TX_DATA_69_const_net_10;
wire   [3:0]     TX_DATA_70_const_net_10;
wire   [3:0]     TX_DATA_71_const_net_10;
wire   [3:0]     TX_DATA_72_const_net_10;
wire   [3:0]     TX_DATA_73_const_net_10;
wire   [3:0]     TX_DATA_74_const_net_10;
wire   [3:0]     TX_DATA_75_const_net_10;
wire   [3:0]     TX_DATA_76_const_net_10;
wire   [3:0]     TX_DATA_77_const_net_10;
wire   [3:0]     TX_DATA_78_const_net_10;
wire   [3:0]     TX_DATA_79_const_net_10;
wire   [3:0]     TX_DATA_80_const_net_10;
wire   [3:0]     TX_DATA_81_const_net_10;
wire   [3:0]     TX_DATA_82_const_net_10;
wire   [3:0]     TX_DATA_83_const_net_10;
wire   [3:0]     TX_DATA_84_const_net_10;
wire   [3:0]     TX_DATA_85_const_net_10;
wire   [3:0]     TX_DATA_86_const_net_10;
wire   [3:0]     TX_DATA_87_const_net_10;
wire   [3:0]     TX_DATA_88_const_net_10;
wire   [3:0]     TX_DATA_89_const_net_10;
wire   [3:0]     TX_DATA_90_const_net_10;
wire   [3:0]     TX_DATA_91_const_net_10;
wire   [3:0]     TX_DATA_92_const_net_10;
wire   [3:0]     TX_DATA_93_const_net_10;
wire   [3:0]     TX_DATA_94_const_net_10;
wire   [3:0]     TX_DATA_95_const_net_10;
wire   [3:0]     TX_DATA_96_const_net_10;
wire   [3:0]     TX_DATA_97_const_net_10;
wire   [3:0]     TX_DATA_98_const_net_10;
wire   [3:0]     TX_DATA_99_const_net_10;
wire   [3:0]     TX_DATA_100_const_net_10;
wire   [3:0]     TX_DATA_101_const_net_10;
wire   [3:0]     TX_DATA_102_const_net_10;
wire   [3:0]     TX_DATA_103_const_net_10;
wire   [3:0]     TX_DATA_104_const_net_10;
wire   [3:0]     TX_DATA_105_const_net_10;
wire   [3:0]     TX_DATA_106_const_net_10;
wire   [3:0]     TX_DATA_107_const_net_10;
wire   [3:0]     TX_DATA_108_const_net_10;
wire   [3:0]     TX_DATA_109_const_net_10;
wire   [3:0]     TX_DATA_110_const_net_10;
wire   [3:0]     TX_DATA_111_const_net_10;
wire   [3:0]     TX_DATA_112_const_net_10;
wire   [3:0]     TX_DATA_113_const_net_10;
wire   [3:0]     TX_DATA_114_const_net_10;
wire   [3:0]     TX_DATA_115_const_net_10;
wire   [3:0]     TX_DATA_116_const_net_10;
wire   [3:0]     TX_DATA_117_const_net_10;
wire   [3:0]     TX_DATA_118_const_net_10;
wire   [3:0]     TX_DATA_119_const_net_10;
wire   [3:0]     TX_DATA_120_const_net_10;
wire   [3:0]     TX_DATA_121_const_net_10;
wire   [3:0]     TX_DATA_122_const_net_10;
wire   [3:0]     TX_DATA_123_const_net_10;
wire   [3:0]     TX_DATA_124_const_net_10;
wire   [3:0]     TX_DATA_125_const_net_10;
wire   [3:0]     TX_DATA_126_const_net_10;
wire   [3:0]     TX_DATA_127_const_net_10;
wire   [3:0]     OE_DATA_1_const_net_10;
wire   [3:0]     OE_DATA_2_const_net_10;
wire   [3:0]     OE_DATA_3_const_net_10;
wire   [3:0]     OE_DATA_4_const_net_10;
wire   [3:0]     OE_DATA_5_const_net_10;
wire   [3:0]     OE_DATA_6_const_net_10;
wire   [3:0]     OE_DATA_7_const_net_10;
wire   [3:0]     OE_DATA_8_const_net_10;
wire   [3:0]     OE_DATA_9_const_net_10;
wire   [3:0]     OE_DATA_10_const_net_10;
wire   [3:0]     OE_DATA_11_const_net_10;
wire   [3:0]     OE_DATA_12_const_net_10;
wire   [3:0]     OE_DATA_13_const_net_10;
wire   [3:0]     OE_DATA_14_const_net_10;
wire   [3:0]     OE_DATA_15_const_net_10;
wire   [3:0]     OE_DATA_16_const_net_10;
wire   [3:0]     OE_DATA_17_const_net_10;
wire   [3:0]     OE_DATA_18_const_net_10;
wire   [3:0]     OE_DATA_19_const_net_10;
wire   [3:0]     OE_DATA_20_const_net_10;
wire   [3:0]     OE_DATA_21_const_net_10;
wire   [3:0]     OE_DATA_22_const_net_10;
wire   [3:0]     OE_DATA_23_const_net_10;
wire   [3:0]     OE_DATA_24_const_net_10;
wire   [3:0]     OE_DATA_25_const_net_10;
wire   [3:0]     OE_DATA_26_const_net_10;
wire   [3:0]     OE_DATA_27_const_net_10;
wire   [3:0]     OE_DATA_28_const_net_10;
wire   [3:0]     OE_DATA_29_const_net_10;
wire   [3:0]     OE_DATA_30_const_net_10;
wire   [3:0]     OE_DATA_31_const_net_10;
wire   [3:0]     OE_DATA_32_const_net_10;
wire   [3:0]     OE_DATA_33_const_net_10;
wire   [3:0]     OE_DATA_34_const_net_10;
wire   [3:0]     OE_DATA_35_const_net_10;
wire   [3:0]     OE_DATA_36_const_net_10;
wire   [3:0]     OE_DATA_37_const_net_10;
wire   [3:0]     OE_DATA_38_const_net_10;
wire   [3:0]     OE_DATA_39_const_net_10;
wire   [3:0]     OE_DATA_40_const_net_10;
wire   [3:0]     OE_DATA_41_const_net_10;
wire   [3:0]     OE_DATA_42_const_net_10;
wire   [3:0]     OE_DATA_43_const_net_10;
wire   [3:0]     OE_DATA_44_const_net_10;
wire   [3:0]     OE_DATA_45_const_net_10;
wire   [3:0]     OE_DATA_46_const_net_10;
wire   [3:0]     OE_DATA_47_const_net_10;
wire   [3:0]     OE_DATA_48_const_net_10;
wire   [3:0]     OE_DATA_49_const_net_10;
wire   [3:0]     OE_DATA_50_const_net_10;
wire   [3:0]     OE_DATA_51_const_net_10;
wire   [3:0]     OE_DATA_52_const_net_10;
wire   [3:0]     OE_DATA_53_const_net_10;
wire   [3:0]     OE_DATA_54_const_net_10;
wire   [3:0]     OE_DATA_55_const_net_10;
wire   [3:0]     OE_DATA_56_const_net_10;
wire   [3:0]     OE_DATA_57_const_net_10;
wire   [3:0]     OE_DATA_58_const_net_10;
wire   [3:0]     OE_DATA_59_const_net_10;
wire   [3:0]     OE_DATA_60_const_net_10;
wire   [3:0]     OE_DATA_61_const_net_10;
wire   [3:0]     OE_DATA_62_const_net_10;
wire   [3:0]     OE_DATA_63_const_net_10;
wire   [3:0]     OE_DATA_64_const_net_10;
wire   [3:0]     OE_DATA_65_const_net_10;
wire   [3:0]     OE_DATA_66_const_net_10;
wire   [3:0]     OE_DATA_67_const_net_10;
wire   [3:0]     OE_DATA_68_const_net_10;
wire   [3:0]     OE_DATA_69_const_net_10;
wire   [3:0]     OE_DATA_70_const_net_10;
wire   [3:0]     OE_DATA_71_const_net_10;
wire   [3:0]     OE_DATA_72_const_net_10;
wire   [3:0]     OE_DATA_73_const_net_10;
wire   [3:0]     OE_DATA_74_const_net_10;
wire   [3:0]     OE_DATA_75_const_net_10;
wire   [3:0]     OE_DATA_76_const_net_10;
wire   [3:0]     OE_DATA_77_const_net_10;
wire   [3:0]     OE_DATA_78_const_net_10;
wire   [3:0]     OE_DATA_79_const_net_10;
wire   [3:0]     OE_DATA_80_const_net_10;
wire   [3:0]     OE_DATA_81_const_net_10;
wire   [3:0]     OE_DATA_82_const_net_10;
wire   [3:0]     OE_DATA_83_const_net_10;
wire   [3:0]     OE_DATA_84_const_net_10;
wire   [3:0]     OE_DATA_85_const_net_10;
wire   [3:0]     OE_DATA_86_const_net_10;
wire   [3:0]     OE_DATA_87_const_net_10;
wire   [3:0]     OE_DATA_88_const_net_10;
wire   [3:0]     OE_DATA_89_const_net_10;
wire   [3:0]     OE_DATA_90_const_net_10;
wire   [3:0]     OE_DATA_91_const_net_10;
wire   [3:0]     OE_DATA_92_const_net_10;
wire   [3:0]     OE_DATA_93_const_net_10;
wire   [3:0]     OE_DATA_94_const_net_10;
wire   [3:0]     OE_DATA_95_const_net_10;
wire   [3:0]     OE_DATA_96_const_net_10;
wire   [3:0]     OE_DATA_97_const_net_10;
wire   [3:0]     OE_DATA_98_const_net_10;
wire   [3:0]     OE_DATA_99_const_net_10;
wire   [3:0]     OE_DATA_100_const_net_10;
wire   [3:0]     OE_DATA_101_const_net_10;
wire   [3:0]     OE_DATA_102_const_net_10;
wire   [3:0]     OE_DATA_103_const_net_10;
wire   [3:0]     OE_DATA_104_const_net_10;
wire   [3:0]     OE_DATA_105_const_net_10;
wire   [3:0]     OE_DATA_106_const_net_10;
wire   [3:0]     OE_DATA_107_const_net_10;
wire   [3:0]     OE_DATA_108_const_net_10;
wire   [3:0]     OE_DATA_109_const_net_10;
wire   [3:0]     OE_DATA_110_const_net_10;
wire   [3:0]     OE_DATA_111_const_net_10;
wire   [3:0]     OE_DATA_112_const_net_10;
wire   [3:0]     OE_DATA_113_const_net_10;
wire   [3:0]     OE_DATA_114_const_net_10;
wire   [3:0]     OE_DATA_115_const_net_10;
wire   [3:0]     OE_DATA_116_const_net_10;
wire   [3:0]     OE_DATA_117_const_net_10;
wire   [3:0]     OE_DATA_118_const_net_10;
wire   [3:0]     OE_DATA_119_const_net_10;
wire   [3:0]     OE_DATA_120_const_net_10;
wire   [3:0]     OE_DATA_121_const_net_10;
wire   [3:0]     OE_DATA_122_const_net_10;
wire   [3:0]     OE_DATA_123_const_net_10;
wire   [3:0]     OE_DATA_124_const_net_10;
wire   [3:0]     OE_DATA_125_const_net_10;
wire   [3:0]     OE_DATA_126_const_net_10;
wire   [3:0]     OE_DATA_127_const_net_10;
wire   [1:0]     RX_DQS_90_const_net_11;
wire   [2:0]     FIFO_WR_PTR_const_net_11;
wire   [2:0]     FIFO_RD_PTR_const_net_11;
wire   [2:0]     EYE_MONITOR_LANE_WIDTH_const_net_11;
wire   [3:0]     TX_DATA_1_const_net_8;
wire   [3:0]     TX_DATA_2_const_net_10;
wire   [3:0]     TX_DATA_3_const_net_10;
wire   [3:0]     TX_DATA_4_const_net_10;
wire   [3:0]     TX_DATA_5_const_net_10;
wire   [3:0]     TX_DATA_6_const_net_10;
wire   [3:0]     TX_DATA_7_const_net_10;
wire   [3:0]     TX_DATA_8_const_net_10;
wire   [3:0]     TX_DATA_9_const_net_10;
wire   [3:0]     TX_DATA_10_const_net_10;
wire   [3:0]     TX_DATA_11_const_net_10;
wire   [3:0]     TX_DATA_12_const_net_11;
wire   [3:0]     TX_DATA_13_const_net_11;
wire   [3:0]     TX_DATA_14_const_net_11;
wire   [3:0]     TX_DATA_15_const_net_11;
wire   [3:0]     TX_DATA_16_const_net_11;
wire   [3:0]     TX_DATA_17_const_net_11;
wire   [3:0]     TX_DATA_18_const_net_11;
wire   [3:0]     TX_DATA_19_const_net_11;
wire   [3:0]     TX_DATA_20_const_net_11;
wire   [3:0]     TX_DATA_21_const_net_11;
wire   [3:0]     TX_DATA_22_const_net_11;
wire   [3:0]     TX_DATA_23_const_net_11;
wire   [3:0]     TX_DATA_24_const_net_11;
wire   [3:0]     TX_DATA_25_const_net_11;
wire   [3:0]     TX_DATA_26_const_net_11;
wire   [3:0]     TX_DATA_27_const_net_11;
wire   [3:0]     TX_DATA_28_const_net_11;
wire   [3:0]     TX_DATA_29_const_net_11;
wire   [3:0]     TX_DATA_30_const_net_11;
wire   [3:0]     TX_DATA_31_const_net_11;
wire   [3:0]     TX_DATA_32_const_net_11;
wire   [3:0]     TX_DATA_33_const_net_11;
wire   [3:0]     TX_DATA_34_const_net_11;
wire   [3:0]     TX_DATA_35_const_net_11;
wire   [3:0]     TX_DATA_36_const_net_11;
wire   [3:0]     TX_DATA_37_const_net_11;
wire   [3:0]     TX_DATA_38_const_net_11;
wire   [3:0]     TX_DATA_39_const_net_11;
wire   [3:0]     TX_DATA_40_const_net_11;
wire   [3:0]     TX_DATA_41_const_net_11;
wire   [3:0]     TX_DATA_42_const_net_11;
wire   [3:0]     TX_DATA_43_const_net_11;
wire   [3:0]     TX_DATA_44_const_net_11;
wire   [3:0]     TX_DATA_45_const_net_11;
wire   [3:0]     TX_DATA_46_const_net_11;
wire   [3:0]     TX_DATA_47_const_net_11;
wire   [3:0]     TX_DATA_48_const_net_11;
wire   [3:0]     TX_DATA_49_const_net_11;
wire   [3:0]     TX_DATA_50_const_net_11;
wire   [3:0]     TX_DATA_51_const_net_11;
wire   [3:0]     TX_DATA_52_const_net_11;
wire   [3:0]     TX_DATA_53_const_net_11;
wire   [3:0]     TX_DATA_54_const_net_11;
wire   [3:0]     TX_DATA_55_const_net_11;
wire   [3:0]     TX_DATA_56_const_net_11;
wire   [3:0]     TX_DATA_57_const_net_11;
wire   [3:0]     TX_DATA_58_const_net_11;
wire   [3:0]     TX_DATA_59_const_net_11;
wire   [3:0]     TX_DATA_60_const_net_11;
wire   [3:0]     TX_DATA_61_const_net_11;
wire   [3:0]     TX_DATA_62_const_net_11;
wire   [3:0]     TX_DATA_63_const_net_11;
wire   [3:0]     TX_DATA_64_const_net_11;
wire   [3:0]     TX_DATA_65_const_net_11;
wire   [3:0]     TX_DATA_66_const_net_11;
wire   [3:0]     TX_DATA_67_const_net_11;
wire   [3:0]     TX_DATA_68_const_net_11;
wire   [3:0]     TX_DATA_69_const_net_11;
wire   [3:0]     TX_DATA_70_const_net_11;
wire   [3:0]     TX_DATA_71_const_net_11;
wire   [3:0]     TX_DATA_72_const_net_11;
wire   [3:0]     TX_DATA_73_const_net_11;
wire   [3:0]     TX_DATA_74_const_net_11;
wire   [3:0]     TX_DATA_75_const_net_11;
wire   [3:0]     TX_DATA_76_const_net_11;
wire   [3:0]     TX_DATA_77_const_net_11;
wire   [3:0]     TX_DATA_78_const_net_11;
wire   [3:0]     TX_DATA_79_const_net_11;
wire   [3:0]     TX_DATA_80_const_net_11;
wire   [3:0]     TX_DATA_81_const_net_11;
wire   [3:0]     TX_DATA_82_const_net_11;
wire   [3:0]     TX_DATA_83_const_net_11;
wire   [3:0]     TX_DATA_84_const_net_11;
wire   [3:0]     TX_DATA_85_const_net_11;
wire   [3:0]     TX_DATA_86_const_net_11;
wire   [3:0]     TX_DATA_87_const_net_11;
wire   [3:0]     TX_DATA_88_const_net_11;
wire   [3:0]     TX_DATA_89_const_net_11;
wire   [3:0]     TX_DATA_90_const_net_11;
wire   [3:0]     TX_DATA_91_const_net_11;
wire   [3:0]     TX_DATA_92_const_net_11;
wire   [3:0]     TX_DATA_93_const_net_11;
wire   [3:0]     TX_DATA_94_const_net_11;
wire   [3:0]     TX_DATA_95_const_net_11;
wire   [3:0]     TX_DATA_96_const_net_11;
wire   [3:0]     TX_DATA_97_const_net_11;
wire   [3:0]     TX_DATA_98_const_net_11;
wire   [3:0]     TX_DATA_99_const_net_11;
wire   [3:0]     TX_DATA_100_const_net_11;
wire   [3:0]     TX_DATA_101_const_net_11;
wire   [3:0]     TX_DATA_102_const_net_11;
wire   [3:0]     TX_DATA_103_const_net_11;
wire   [3:0]     TX_DATA_104_const_net_11;
wire   [3:0]     TX_DATA_105_const_net_11;
wire   [3:0]     TX_DATA_106_const_net_11;
wire   [3:0]     TX_DATA_107_const_net_11;
wire   [3:0]     TX_DATA_108_const_net_11;
wire   [3:0]     TX_DATA_109_const_net_11;
wire   [3:0]     TX_DATA_110_const_net_11;
wire   [3:0]     TX_DATA_111_const_net_11;
wire   [3:0]     TX_DATA_112_const_net_11;
wire   [3:0]     TX_DATA_113_const_net_11;
wire   [3:0]     TX_DATA_114_const_net_11;
wire   [3:0]     TX_DATA_115_const_net_11;
wire   [3:0]     TX_DATA_116_const_net_11;
wire   [3:0]     TX_DATA_117_const_net_11;
wire   [3:0]     TX_DATA_118_const_net_11;
wire   [3:0]     TX_DATA_119_const_net_11;
wire   [3:0]     TX_DATA_120_const_net_11;
wire   [3:0]     TX_DATA_121_const_net_11;
wire   [3:0]     TX_DATA_122_const_net_11;
wire   [3:0]     TX_DATA_123_const_net_11;
wire   [3:0]     TX_DATA_124_const_net_11;
wire   [3:0]     TX_DATA_125_const_net_11;
wire   [3:0]     TX_DATA_126_const_net_11;
wire   [3:0]     TX_DATA_127_const_net_11;
wire   [3:0]     OE_DATA_1_const_net_11;
wire   [3:0]     OE_DATA_2_const_net_11;
wire   [3:0]     OE_DATA_3_const_net_11;
wire   [3:0]     OE_DATA_4_const_net_11;
wire   [3:0]     OE_DATA_5_const_net_11;
wire   [3:0]     OE_DATA_6_const_net_11;
wire   [3:0]     OE_DATA_7_const_net_11;
wire   [3:0]     OE_DATA_8_const_net_11;
wire   [3:0]     OE_DATA_9_const_net_11;
wire   [3:0]     OE_DATA_10_const_net_11;
wire   [3:0]     OE_DATA_11_const_net_11;
wire   [3:0]     OE_DATA_12_const_net_11;
wire   [3:0]     OE_DATA_13_const_net_11;
wire   [3:0]     OE_DATA_14_const_net_11;
wire   [3:0]     OE_DATA_15_const_net_11;
wire   [3:0]     OE_DATA_16_const_net_11;
wire   [3:0]     OE_DATA_17_const_net_11;
wire   [3:0]     OE_DATA_18_const_net_11;
wire   [3:0]     OE_DATA_19_const_net_11;
wire   [3:0]     OE_DATA_20_const_net_11;
wire   [3:0]     OE_DATA_21_const_net_11;
wire   [3:0]     OE_DATA_22_const_net_11;
wire   [3:0]     OE_DATA_23_const_net_11;
wire   [3:0]     OE_DATA_24_const_net_11;
wire   [3:0]     OE_DATA_25_const_net_11;
wire   [3:0]     OE_DATA_26_const_net_11;
wire   [3:0]     OE_DATA_27_const_net_11;
wire   [3:0]     OE_DATA_28_const_net_11;
wire   [3:0]     OE_DATA_29_const_net_11;
wire   [3:0]     OE_DATA_30_const_net_11;
wire   [3:0]     OE_DATA_31_const_net_11;
wire   [3:0]     OE_DATA_32_const_net_11;
wire   [3:0]     OE_DATA_33_const_net_11;
wire   [3:0]     OE_DATA_34_const_net_11;
wire   [3:0]     OE_DATA_35_const_net_11;
wire   [3:0]     OE_DATA_36_const_net_11;
wire   [3:0]     OE_DATA_37_const_net_11;
wire   [3:0]     OE_DATA_38_const_net_11;
wire   [3:0]     OE_DATA_39_const_net_11;
wire   [3:0]     OE_DATA_40_const_net_11;
wire   [3:0]     OE_DATA_41_const_net_11;
wire   [3:0]     OE_DATA_42_const_net_11;
wire   [3:0]     OE_DATA_43_const_net_11;
wire   [3:0]     OE_DATA_44_const_net_11;
wire   [3:0]     OE_DATA_45_const_net_11;
wire   [3:0]     OE_DATA_46_const_net_11;
wire   [3:0]     OE_DATA_47_const_net_11;
wire   [3:0]     OE_DATA_48_const_net_11;
wire   [3:0]     OE_DATA_49_const_net_11;
wire   [3:0]     OE_DATA_50_const_net_11;
wire   [3:0]     OE_DATA_51_const_net_11;
wire   [3:0]     OE_DATA_52_const_net_11;
wire   [3:0]     OE_DATA_53_const_net_11;
wire   [3:0]     OE_DATA_54_const_net_11;
wire   [3:0]     OE_DATA_55_const_net_11;
wire   [3:0]     OE_DATA_56_const_net_11;
wire   [3:0]     OE_DATA_57_const_net_11;
wire   [3:0]     OE_DATA_58_const_net_11;
wire   [3:0]     OE_DATA_59_const_net_11;
wire   [3:0]     OE_DATA_60_const_net_11;
wire   [3:0]     OE_DATA_61_const_net_11;
wire   [3:0]     OE_DATA_62_const_net_11;
wire   [3:0]     OE_DATA_63_const_net_11;
wire   [3:0]     OE_DATA_64_const_net_11;
wire   [3:0]     OE_DATA_65_const_net_11;
wire   [3:0]     OE_DATA_66_const_net_11;
wire   [3:0]     OE_DATA_67_const_net_11;
wire   [3:0]     OE_DATA_68_const_net_11;
wire   [3:0]     OE_DATA_69_const_net_11;
wire   [3:0]     OE_DATA_70_const_net_11;
wire   [3:0]     OE_DATA_71_const_net_11;
wire   [3:0]     OE_DATA_72_const_net_11;
wire   [3:0]     OE_DATA_73_const_net_11;
wire   [3:0]     OE_DATA_74_const_net_11;
wire   [3:0]     OE_DATA_75_const_net_11;
wire   [3:0]     OE_DATA_76_const_net_11;
wire   [3:0]     OE_DATA_77_const_net_11;
wire   [3:0]     OE_DATA_78_const_net_11;
wire   [3:0]     OE_DATA_79_const_net_11;
wire   [3:0]     OE_DATA_80_const_net_11;
wire   [3:0]     OE_DATA_81_const_net_11;
wire   [3:0]     OE_DATA_82_const_net_11;
wire   [3:0]     OE_DATA_83_const_net_11;
wire   [3:0]     OE_DATA_84_const_net_11;
wire   [3:0]     OE_DATA_85_const_net_11;
wire   [3:0]     OE_DATA_86_const_net_11;
wire   [3:0]     OE_DATA_87_const_net_11;
wire   [3:0]     OE_DATA_88_const_net_11;
wire   [3:0]     OE_DATA_89_const_net_11;
wire   [3:0]     OE_DATA_90_const_net_11;
wire   [3:0]     OE_DATA_91_const_net_11;
wire   [3:0]     OE_DATA_92_const_net_11;
wire   [3:0]     OE_DATA_93_const_net_11;
wire   [3:0]     OE_DATA_94_const_net_11;
wire   [3:0]     OE_DATA_95_const_net_11;
wire   [3:0]     OE_DATA_96_const_net_11;
wire   [3:0]     OE_DATA_97_const_net_11;
wire   [3:0]     OE_DATA_98_const_net_11;
wire   [3:0]     OE_DATA_99_const_net_11;
wire   [3:0]     OE_DATA_100_const_net_11;
wire   [3:0]     OE_DATA_101_const_net_11;
wire   [3:0]     OE_DATA_102_const_net_11;
wire   [3:0]     OE_DATA_103_const_net_11;
wire   [3:0]     OE_DATA_104_const_net_11;
wire   [3:0]     OE_DATA_105_const_net_11;
wire   [3:0]     OE_DATA_106_const_net_11;
wire   [3:0]     OE_DATA_107_const_net_11;
wire   [3:0]     OE_DATA_108_const_net_11;
wire   [3:0]     OE_DATA_109_const_net_11;
wire   [3:0]     OE_DATA_110_const_net_11;
wire   [3:0]     OE_DATA_111_const_net_11;
wire   [3:0]     OE_DATA_112_const_net_11;
wire   [3:0]     OE_DATA_113_const_net_11;
wire   [3:0]     OE_DATA_114_const_net_11;
wire   [3:0]     OE_DATA_115_const_net_11;
wire   [3:0]     OE_DATA_116_const_net_11;
wire   [3:0]     OE_DATA_117_const_net_11;
wire   [3:0]     OE_DATA_118_const_net_11;
wire   [3:0]     OE_DATA_119_const_net_11;
wire   [3:0]     OE_DATA_120_const_net_11;
wire   [3:0]     OE_DATA_121_const_net_11;
wire   [3:0]     OE_DATA_122_const_net_11;
wire   [3:0]     OE_DATA_123_const_net_11;
wire   [3:0]     OE_DATA_124_const_net_11;
wire   [3:0]     OE_DATA_125_const_net_11;
wire   [3:0]     OE_DATA_126_const_net_11;
wire   [3:0]     OE_DATA_127_const_net_11;
wire   [1:0]     RX_DQS_90_const_net_12;
wire   [2:0]     FIFO_WR_PTR_const_net_12;
wire   [2:0]     FIFO_RD_PTR_const_net_12;
wire   [2:0]     EYE_MONITOR_LANE_WIDTH_const_net_12;
wire   [7:0]     TX_DATA_0_const_net_9;
wire   [7:0]     TX_DATA_1_const_net_9;
wire   [7:0]     TX_DATA_2_const_net_11;
wire   [7:0]     TX_DATA_3_const_net_11;
wire   [7:0]     TX_DATA_4_const_net_11;
wire   [7:0]     TX_DATA_5_const_net_11;
wire   [7:0]     TX_DATA_6_const_net_11;
wire   [7:0]     TX_DATA_7_const_net_11;
wire   [7:0]     TX_DATA_8_const_net_11;
wire   [7:0]     TX_DATA_9_const_net_11;
wire   [7:0]     TX_DATA_10_const_net_11;
wire   [7:0]     TX_DATA_11_const_net_11;
wire   [7:0]     TX_DATA_12_const_net_12;
wire   [7:0]     TX_DATA_13_const_net_12;
wire   [7:0]     TX_DATA_14_const_net_12;
wire   [7:0]     TX_DATA_15_const_net_12;
wire   [7:0]     TX_DATA_16_const_net_12;
wire   [7:0]     TX_DATA_17_const_net_12;
wire   [7:0]     TX_DATA_18_const_net_12;
wire   [7:0]     TX_DATA_19_const_net_12;
wire   [7:0]     TX_DATA_20_const_net_12;
wire   [7:0]     TX_DATA_21_const_net_12;
wire   [7:0]     TX_DATA_22_const_net_12;
wire   [7:0]     TX_DATA_23_const_net_12;
wire   [7:0]     TX_DATA_24_const_net_12;
wire   [7:0]     TX_DATA_25_const_net_12;
wire   [7:0]     TX_DATA_26_const_net_12;
wire   [7:0]     TX_DATA_27_const_net_12;
wire   [7:0]     TX_DATA_28_const_net_12;
wire   [7:0]     TX_DATA_29_const_net_12;
wire   [7:0]     TX_DATA_30_const_net_12;
wire   [7:0]     TX_DATA_31_const_net_12;
wire   [7:0]     TX_DATA_32_const_net_12;
wire   [7:0]     TX_DATA_33_const_net_12;
wire   [7:0]     TX_DATA_34_const_net_12;
wire   [7:0]     TX_DATA_35_const_net_12;
wire   [7:0]     TX_DATA_36_const_net_12;
wire   [7:0]     TX_DATA_37_const_net_12;
wire   [7:0]     TX_DATA_38_const_net_12;
wire   [7:0]     TX_DATA_39_const_net_12;
wire   [7:0]     TX_DATA_40_const_net_12;
wire   [7:0]     TX_DATA_41_const_net_12;
wire   [7:0]     TX_DATA_42_const_net_12;
wire   [7:0]     TX_DATA_43_const_net_12;
wire   [7:0]     TX_DATA_44_const_net_12;
wire   [7:0]     TX_DATA_45_const_net_12;
wire   [7:0]     TX_DATA_46_const_net_12;
wire   [7:0]     TX_DATA_47_const_net_12;
wire   [7:0]     TX_DATA_48_const_net_12;
wire   [7:0]     TX_DATA_49_const_net_12;
wire   [7:0]     TX_DATA_50_const_net_12;
wire   [7:0]     TX_DATA_51_const_net_12;
wire   [7:0]     TX_DATA_52_const_net_12;
wire   [7:0]     TX_DATA_53_const_net_12;
wire   [7:0]     TX_DATA_54_const_net_12;
wire   [7:0]     TX_DATA_55_const_net_12;
wire   [7:0]     TX_DATA_56_const_net_12;
wire   [7:0]     TX_DATA_57_const_net_12;
wire   [7:0]     TX_DATA_58_const_net_12;
wire   [7:0]     TX_DATA_59_const_net_12;
wire   [7:0]     TX_DATA_60_const_net_12;
wire   [7:0]     TX_DATA_61_const_net_12;
wire   [7:0]     TX_DATA_62_const_net_12;
wire   [7:0]     TX_DATA_63_const_net_12;
wire   [7:0]     TX_DATA_64_const_net_12;
wire   [7:0]     TX_DATA_65_const_net_12;
wire   [7:0]     TX_DATA_66_const_net_12;
wire   [7:0]     TX_DATA_67_const_net_12;
wire   [7:0]     TX_DATA_68_const_net_12;
wire   [7:0]     TX_DATA_69_const_net_12;
wire   [7:0]     TX_DATA_70_const_net_12;
wire   [7:0]     TX_DATA_71_const_net_12;
wire   [7:0]     TX_DATA_72_const_net_12;
wire   [7:0]     TX_DATA_73_const_net_12;
wire   [7:0]     TX_DATA_74_const_net_12;
wire   [7:0]     TX_DATA_75_const_net_12;
wire   [7:0]     TX_DATA_76_const_net_12;
wire   [7:0]     TX_DATA_77_const_net_12;
wire   [7:0]     TX_DATA_78_const_net_12;
wire   [7:0]     TX_DATA_79_const_net_12;
wire   [7:0]     TX_DATA_80_const_net_12;
wire   [7:0]     TX_DATA_81_const_net_12;
wire   [7:0]     TX_DATA_82_const_net_12;
wire   [7:0]     TX_DATA_83_const_net_12;
wire   [7:0]     TX_DATA_84_const_net_12;
wire   [7:0]     TX_DATA_85_const_net_12;
wire   [7:0]     TX_DATA_86_const_net_12;
wire   [7:0]     TX_DATA_87_const_net_12;
wire   [7:0]     TX_DATA_88_const_net_12;
wire   [7:0]     TX_DATA_89_const_net_12;
wire   [7:0]     TX_DATA_90_const_net_12;
wire   [7:0]     TX_DATA_91_const_net_12;
wire   [7:0]     TX_DATA_92_const_net_12;
wire   [7:0]     TX_DATA_93_const_net_12;
wire   [7:0]     TX_DATA_94_const_net_12;
wire   [7:0]     TX_DATA_95_const_net_12;
wire   [7:0]     TX_DATA_96_const_net_12;
wire   [7:0]     TX_DATA_97_const_net_12;
wire   [7:0]     TX_DATA_98_const_net_12;
wire   [7:0]     TX_DATA_99_const_net_12;
wire   [7:0]     TX_DATA_100_const_net_12;
wire   [7:0]     TX_DATA_101_const_net_12;
wire   [7:0]     TX_DATA_102_const_net_12;
wire   [7:0]     TX_DATA_103_const_net_12;
wire   [7:0]     TX_DATA_104_const_net_12;
wire   [7:0]     TX_DATA_105_const_net_12;
wire   [7:0]     TX_DATA_106_const_net_12;
wire   [7:0]     TX_DATA_107_const_net_12;
wire   [7:0]     TX_DATA_108_const_net_12;
wire   [7:0]     TX_DATA_109_const_net_12;
wire   [7:0]     TX_DATA_110_const_net_12;
wire   [7:0]     TX_DATA_111_const_net_12;
wire   [7:0]     TX_DATA_112_const_net_12;
wire   [7:0]     TX_DATA_113_const_net_12;
wire   [7:0]     TX_DATA_114_const_net_12;
wire   [7:0]     TX_DATA_115_const_net_12;
wire   [7:0]     TX_DATA_116_const_net_12;
wire   [7:0]     TX_DATA_117_const_net_12;
wire   [7:0]     TX_DATA_118_const_net_12;
wire   [7:0]     TX_DATA_119_const_net_12;
wire   [7:0]     TX_DATA_120_const_net_12;
wire   [7:0]     TX_DATA_121_const_net_12;
wire   [7:0]     TX_DATA_122_const_net_12;
wire   [7:0]     TX_DATA_123_const_net_12;
wire   [7:0]     TX_DATA_124_const_net_12;
wire   [7:0]     TX_DATA_125_const_net_12;
wire   [7:0]     TX_DATA_126_const_net_12;
wire   [7:0]     TX_DATA_127_const_net_12;
wire   [3:0]     OE_DATA_0_const_net_17;
wire   [3:0]     OE_DATA_1_const_net_12;
wire   [3:0]     OE_DATA_2_const_net_12;
wire   [3:0]     OE_DATA_3_const_net_12;
wire   [3:0]     OE_DATA_4_const_net_12;
wire   [3:0]     OE_DATA_5_const_net_12;
wire   [3:0]     OE_DATA_6_const_net_12;
wire   [3:0]     OE_DATA_7_const_net_12;
wire   [3:0]     OE_DATA_8_const_net_12;
wire   [3:0]     OE_DATA_9_const_net_12;
wire   [3:0]     OE_DATA_10_const_net_12;
wire   [3:0]     OE_DATA_11_const_net_12;
wire   [3:0]     OE_DATA_12_const_net_12;
wire   [3:0]     OE_DATA_13_const_net_12;
wire   [3:0]     OE_DATA_14_const_net_12;
wire   [3:0]     OE_DATA_15_const_net_12;
wire   [3:0]     OE_DATA_16_const_net_12;
wire   [3:0]     OE_DATA_17_const_net_12;
wire   [3:0]     OE_DATA_18_const_net_12;
wire   [3:0]     OE_DATA_19_const_net_12;
wire   [3:0]     OE_DATA_20_const_net_12;
wire   [3:0]     OE_DATA_21_const_net_12;
wire   [3:0]     OE_DATA_22_const_net_12;
wire   [3:0]     OE_DATA_23_const_net_12;
wire   [3:0]     OE_DATA_24_const_net_12;
wire   [3:0]     OE_DATA_25_const_net_12;
wire   [3:0]     OE_DATA_26_const_net_12;
wire   [3:0]     OE_DATA_27_const_net_12;
wire   [3:0]     OE_DATA_28_const_net_12;
wire   [3:0]     OE_DATA_29_const_net_12;
wire   [3:0]     OE_DATA_30_const_net_12;
wire   [3:0]     OE_DATA_31_const_net_12;
wire   [3:0]     OE_DATA_32_const_net_12;
wire   [3:0]     OE_DATA_33_const_net_12;
wire   [3:0]     OE_DATA_34_const_net_12;
wire   [3:0]     OE_DATA_35_const_net_12;
wire   [3:0]     OE_DATA_36_const_net_12;
wire   [3:0]     OE_DATA_37_const_net_12;
wire   [3:0]     OE_DATA_38_const_net_12;
wire   [3:0]     OE_DATA_39_const_net_12;
wire   [3:0]     OE_DATA_40_const_net_12;
wire   [3:0]     OE_DATA_41_const_net_12;
wire   [3:0]     OE_DATA_42_const_net_12;
wire   [3:0]     OE_DATA_43_const_net_12;
wire   [3:0]     OE_DATA_44_const_net_12;
wire   [3:0]     OE_DATA_45_const_net_12;
wire   [3:0]     OE_DATA_46_const_net_12;
wire   [3:0]     OE_DATA_47_const_net_12;
wire   [3:0]     OE_DATA_48_const_net_12;
wire   [3:0]     OE_DATA_49_const_net_12;
wire   [3:0]     OE_DATA_50_const_net_12;
wire   [3:0]     OE_DATA_51_const_net_12;
wire   [3:0]     OE_DATA_52_const_net_12;
wire   [3:0]     OE_DATA_53_const_net_12;
wire   [3:0]     OE_DATA_54_const_net_12;
wire   [3:0]     OE_DATA_55_const_net_12;
wire   [3:0]     OE_DATA_56_const_net_12;
wire   [3:0]     OE_DATA_57_const_net_12;
wire   [3:0]     OE_DATA_58_const_net_12;
wire   [3:0]     OE_DATA_59_const_net_12;
wire   [3:0]     OE_DATA_60_const_net_12;
wire   [3:0]     OE_DATA_61_const_net_12;
wire   [3:0]     OE_DATA_62_const_net_12;
wire   [3:0]     OE_DATA_63_const_net_12;
wire   [3:0]     OE_DATA_64_const_net_12;
wire   [3:0]     OE_DATA_65_const_net_12;
wire   [3:0]     OE_DATA_66_const_net_12;
wire   [3:0]     OE_DATA_67_const_net_12;
wire   [3:0]     OE_DATA_68_const_net_12;
wire   [3:0]     OE_DATA_69_const_net_12;
wire   [3:0]     OE_DATA_70_const_net_12;
wire   [3:0]     OE_DATA_71_const_net_12;
wire   [3:0]     OE_DATA_72_const_net_12;
wire   [3:0]     OE_DATA_73_const_net_12;
wire   [3:0]     OE_DATA_74_const_net_12;
wire   [3:0]     OE_DATA_75_const_net_12;
wire   [3:0]     OE_DATA_76_const_net_12;
wire   [3:0]     OE_DATA_77_const_net_12;
wire   [3:0]     OE_DATA_78_const_net_12;
wire   [3:0]     OE_DATA_79_const_net_12;
wire   [3:0]     OE_DATA_80_const_net_12;
wire   [3:0]     OE_DATA_81_const_net_12;
wire   [3:0]     OE_DATA_82_const_net_12;
wire   [3:0]     OE_DATA_83_const_net_12;
wire   [3:0]     OE_DATA_84_const_net_12;
wire   [3:0]     OE_DATA_85_const_net_12;
wire   [3:0]     OE_DATA_86_const_net_12;
wire   [3:0]     OE_DATA_87_const_net_12;
wire   [3:0]     OE_DATA_88_const_net_12;
wire   [3:0]     OE_DATA_89_const_net_12;
wire   [3:0]     OE_DATA_90_const_net_12;
wire   [3:0]     OE_DATA_91_const_net_12;
wire   [3:0]     OE_DATA_92_const_net_12;
wire   [3:0]     OE_DATA_93_const_net_12;
wire   [3:0]     OE_DATA_94_const_net_12;
wire   [3:0]     OE_DATA_95_const_net_12;
wire   [3:0]     OE_DATA_96_const_net_12;
wire   [3:0]     OE_DATA_97_const_net_12;
wire   [3:0]     OE_DATA_98_const_net_12;
wire   [3:0]     OE_DATA_99_const_net_12;
wire   [3:0]     OE_DATA_100_const_net_12;
wire   [3:0]     OE_DATA_101_const_net_12;
wire   [3:0]     OE_DATA_102_const_net_12;
wire   [3:0]     OE_DATA_103_const_net_12;
wire   [3:0]     OE_DATA_104_const_net_12;
wire   [3:0]     OE_DATA_105_const_net_12;
wire   [3:0]     OE_DATA_106_const_net_12;
wire   [3:0]     OE_DATA_107_const_net_12;
wire   [3:0]     OE_DATA_108_const_net_12;
wire   [3:0]     OE_DATA_109_const_net_12;
wire   [3:0]     OE_DATA_110_const_net_12;
wire   [3:0]     OE_DATA_111_const_net_12;
wire   [3:0]     OE_DATA_112_const_net_12;
wire   [3:0]     OE_DATA_113_const_net_12;
wire   [3:0]     OE_DATA_114_const_net_12;
wire   [3:0]     OE_DATA_115_const_net_12;
wire   [3:0]     OE_DATA_116_const_net_12;
wire   [3:0]     OE_DATA_117_const_net_12;
wire   [3:0]     OE_DATA_118_const_net_12;
wire   [3:0]     OE_DATA_119_const_net_12;
wire   [3:0]     OE_DATA_120_const_net_12;
wire   [3:0]     OE_DATA_121_const_net_12;
wire   [3:0]     OE_DATA_122_const_net_12;
wire   [3:0]     OE_DATA_123_const_net_12;
wire   [3:0]     OE_DATA_124_const_net_12;
wire   [3:0]     OE_DATA_125_const_net_12;
wire   [3:0]     OE_DATA_126_const_net_12;
wire   [3:0]     OE_DATA_127_const_net_12;
wire   [1:0]     RX_DQS_90_const_net_13;
wire   [2:0]     FIFO_WR_PTR_const_net_13;
wire   [2:0]     FIFO_RD_PTR_const_net_13;
wire   [2:0]     EYE_MONITOR_LANE_WIDTH_const_net_13;
wire   [3:0]     TX_DATA_1_const_net_10;
wire   [3:0]     TX_DATA_2_const_net_12;
wire   [3:0]     TX_DATA_3_const_net_12;
wire   [3:0]     TX_DATA_4_const_net_12;
wire   [3:0]     TX_DATA_5_const_net_12;
wire   [3:0]     TX_DATA_6_const_net_12;
wire   [3:0]     TX_DATA_7_const_net_12;
wire   [3:0]     TX_DATA_8_const_net_12;
wire   [3:0]     TX_DATA_9_const_net_12;
wire   [3:0]     TX_DATA_10_const_net_12;
wire   [3:0]     TX_DATA_11_const_net_12;
wire   [3:0]     TX_DATA_12_const_net_13;
wire   [3:0]     TX_DATA_13_const_net_13;
wire   [3:0]     TX_DATA_14_const_net_13;
wire   [3:0]     TX_DATA_15_const_net_13;
wire   [3:0]     TX_DATA_16_const_net_13;
wire   [3:0]     TX_DATA_17_const_net_13;
wire   [3:0]     TX_DATA_18_const_net_13;
wire   [3:0]     TX_DATA_19_const_net_13;
wire   [3:0]     TX_DATA_20_const_net_13;
wire   [3:0]     TX_DATA_21_const_net_13;
wire   [3:0]     TX_DATA_22_const_net_13;
wire   [3:0]     TX_DATA_23_const_net_13;
wire   [3:0]     TX_DATA_24_const_net_13;
wire   [3:0]     TX_DATA_25_const_net_13;
wire   [3:0]     TX_DATA_26_const_net_13;
wire   [3:0]     TX_DATA_27_const_net_13;
wire   [3:0]     TX_DATA_28_const_net_13;
wire   [3:0]     TX_DATA_29_const_net_13;
wire   [3:0]     TX_DATA_30_const_net_13;
wire   [3:0]     TX_DATA_31_const_net_13;
wire   [3:0]     TX_DATA_32_const_net_13;
wire   [3:0]     TX_DATA_33_const_net_13;
wire   [3:0]     TX_DATA_34_const_net_13;
wire   [3:0]     TX_DATA_35_const_net_13;
wire   [3:0]     TX_DATA_36_const_net_13;
wire   [3:0]     TX_DATA_37_const_net_13;
wire   [3:0]     TX_DATA_38_const_net_13;
wire   [3:0]     TX_DATA_39_const_net_13;
wire   [3:0]     TX_DATA_40_const_net_13;
wire   [3:0]     TX_DATA_41_const_net_13;
wire   [3:0]     TX_DATA_42_const_net_13;
wire   [3:0]     TX_DATA_43_const_net_13;
wire   [3:0]     TX_DATA_44_const_net_13;
wire   [3:0]     TX_DATA_45_const_net_13;
wire   [3:0]     TX_DATA_46_const_net_13;
wire   [3:0]     TX_DATA_47_const_net_13;
wire   [3:0]     TX_DATA_48_const_net_13;
wire   [3:0]     TX_DATA_49_const_net_13;
wire   [3:0]     TX_DATA_50_const_net_13;
wire   [3:0]     TX_DATA_51_const_net_13;
wire   [3:0]     TX_DATA_52_const_net_13;
wire   [3:0]     TX_DATA_53_const_net_13;
wire   [3:0]     TX_DATA_54_const_net_13;
wire   [3:0]     TX_DATA_55_const_net_13;
wire   [3:0]     TX_DATA_56_const_net_13;
wire   [3:0]     TX_DATA_57_const_net_13;
wire   [3:0]     TX_DATA_58_const_net_13;
wire   [3:0]     TX_DATA_59_const_net_13;
wire   [3:0]     TX_DATA_60_const_net_13;
wire   [3:0]     TX_DATA_61_const_net_13;
wire   [3:0]     TX_DATA_62_const_net_13;
wire   [3:0]     TX_DATA_63_const_net_13;
wire   [3:0]     TX_DATA_64_const_net_13;
wire   [3:0]     TX_DATA_65_const_net_13;
wire   [3:0]     TX_DATA_66_const_net_13;
wire   [3:0]     TX_DATA_67_const_net_13;
wire   [3:0]     TX_DATA_68_const_net_13;
wire   [3:0]     TX_DATA_69_const_net_13;
wire   [3:0]     TX_DATA_70_const_net_13;
wire   [3:0]     TX_DATA_71_const_net_13;
wire   [3:0]     TX_DATA_72_const_net_13;
wire   [3:0]     TX_DATA_73_const_net_13;
wire   [3:0]     TX_DATA_74_const_net_13;
wire   [3:0]     TX_DATA_75_const_net_13;
wire   [3:0]     TX_DATA_76_const_net_13;
wire   [3:0]     TX_DATA_77_const_net_13;
wire   [3:0]     TX_DATA_78_const_net_13;
wire   [3:0]     TX_DATA_79_const_net_13;
wire   [3:0]     TX_DATA_80_const_net_13;
wire   [3:0]     TX_DATA_81_const_net_13;
wire   [3:0]     TX_DATA_82_const_net_13;
wire   [3:0]     TX_DATA_83_const_net_13;
wire   [3:0]     TX_DATA_84_const_net_13;
wire   [3:0]     TX_DATA_85_const_net_13;
wire   [3:0]     TX_DATA_86_const_net_13;
wire   [3:0]     TX_DATA_87_const_net_13;
wire   [3:0]     TX_DATA_88_const_net_13;
wire   [3:0]     TX_DATA_89_const_net_13;
wire   [3:0]     TX_DATA_90_const_net_13;
wire   [3:0]     TX_DATA_91_const_net_13;
wire   [3:0]     TX_DATA_92_const_net_13;
wire   [3:0]     TX_DATA_93_const_net_13;
wire   [3:0]     TX_DATA_94_const_net_13;
wire   [3:0]     TX_DATA_95_const_net_13;
wire   [3:0]     TX_DATA_96_const_net_13;
wire   [3:0]     TX_DATA_97_const_net_13;
wire   [3:0]     TX_DATA_98_const_net_13;
wire   [3:0]     TX_DATA_99_const_net_13;
wire   [3:0]     TX_DATA_100_const_net_13;
wire   [3:0]     TX_DATA_101_const_net_13;
wire   [3:0]     TX_DATA_102_const_net_13;
wire   [3:0]     TX_DATA_103_const_net_13;
wire   [3:0]     TX_DATA_104_const_net_13;
wire   [3:0]     TX_DATA_105_const_net_13;
wire   [3:0]     TX_DATA_106_const_net_13;
wire   [3:0]     TX_DATA_107_const_net_13;
wire   [3:0]     TX_DATA_108_const_net_13;
wire   [3:0]     TX_DATA_109_const_net_13;
wire   [3:0]     TX_DATA_110_const_net_13;
wire   [3:0]     TX_DATA_111_const_net_13;
wire   [3:0]     TX_DATA_112_const_net_13;
wire   [3:0]     TX_DATA_113_const_net_13;
wire   [3:0]     TX_DATA_114_const_net_13;
wire   [3:0]     TX_DATA_115_const_net_13;
wire   [3:0]     TX_DATA_116_const_net_13;
wire   [3:0]     TX_DATA_117_const_net_13;
wire   [3:0]     TX_DATA_118_const_net_13;
wire   [3:0]     TX_DATA_119_const_net_13;
wire   [3:0]     TX_DATA_120_const_net_13;
wire   [3:0]     TX_DATA_121_const_net_13;
wire   [3:0]     TX_DATA_122_const_net_13;
wire   [3:0]     TX_DATA_123_const_net_13;
wire   [3:0]     TX_DATA_124_const_net_13;
wire   [3:0]     TX_DATA_125_const_net_13;
wire   [3:0]     TX_DATA_126_const_net_13;
wire   [3:0]     TX_DATA_127_const_net_13;
wire   [3:0]     OE_DATA_1_const_net_13;
wire   [3:0]     OE_DATA_2_const_net_13;
wire   [3:0]     OE_DATA_3_const_net_13;
wire   [3:0]     OE_DATA_4_const_net_13;
wire   [3:0]     OE_DATA_5_const_net_13;
wire   [3:0]     OE_DATA_6_const_net_13;
wire   [3:0]     OE_DATA_7_const_net_13;
wire   [3:0]     OE_DATA_8_const_net_13;
wire   [3:0]     OE_DATA_9_const_net_13;
wire   [3:0]     OE_DATA_10_const_net_13;
wire   [3:0]     OE_DATA_11_const_net_13;
wire   [3:0]     OE_DATA_12_const_net_13;
wire   [3:0]     OE_DATA_13_const_net_13;
wire   [3:0]     OE_DATA_14_const_net_13;
wire   [3:0]     OE_DATA_15_const_net_13;
wire   [3:0]     OE_DATA_16_const_net_13;
wire   [3:0]     OE_DATA_17_const_net_13;
wire   [3:0]     OE_DATA_18_const_net_13;
wire   [3:0]     OE_DATA_19_const_net_13;
wire   [3:0]     OE_DATA_20_const_net_13;
wire   [3:0]     OE_DATA_21_const_net_13;
wire   [3:0]     OE_DATA_22_const_net_13;
wire   [3:0]     OE_DATA_23_const_net_13;
wire   [3:0]     OE_DATA_24_const_net_13;
wire   [3:0]     OE_DATA_25_const_net_13;
wire   [3:0]     OE_DATA_26_const_net_13;
wire   [3:0]     OE_DATA_27_const_net_13;
wire   [3:0]     OE_DATA_28_const_net_13;
wire   [3:0]     OE_DATA_29_const_net_13;
wire   [3:0]     OE_DATA_30_const_net_13;
wire   [3:0]     OE_DATA_31_const_net_13;
wire   [3:0]     OE_DATA_32_const_net_13;
wire   [3:0]     OE_DATA_33_const_net_13;
wire   [3:0]     OE_DATA_34_const_net_13;
wire   [3:0]     OE_DATA_35_const_net_13;
wire   [3:0]     OE_DATA_36_const_net_13;
wire   [3:0]     OE_DATA_37_const_net_13;
wire   [3:0]     OE_DATA_38_const_net_13;
wire   [3:0]     OE_DATA_39_const_net_13;
wire   [3:0]     OE_DATA_40_const_net_13;
wire   [3:0]     OE_DATA_41_const_net_13;
wire   [3:0]     OE_DATA_42_const_net_13;
wire   [3:0]     OE_DATA_43_const_net_13;
wire   [3:0]     OE_DATA_44_const_net_13;
wire   [3:0]     OE_DATA_45_const_net_13;
wire   [3:0]     OE_DATA_46_const_net_13;
wire   [3:0]     OE_DATA_47_const_net_13;
wire   [3:0]     OE_DATA_48_const_net_13;
wire   [3:0]     OE_DATA_49_const_net_13;
wire   [3:0]     OE_DATA_50_const_net_13;
wire   [3:0]     OE_DATA_51_const_net_13;
wire   [3:0]     OE_DATA_52_const_net_13;
wire   [3:0]     OE_DATA_53_const_net_13;
wire   [3:0]     OE_DATA_54_const_net_13;
wire   [3:0]     OE_DATA_55_const_net_13;
wire   [3:0]     OE_DATA_56_const_net_13;
wire   [3:0]     OE_DATA_57_const_net_13;
wire   [3:0]     OE_DATA_58_const_net_13;
wire   [3:0]     OE_DATA_59_const_net_13;
wire   [3:0]     OE_DATA_60_const_net_13;
wire   [3:0]     OE_DATA_61_const_net_13;
wire   [3:0]     OE_DATA_62_const_net_13;
wire   [3:0]     OE_DATA_63_const_net_13;
wire   [3:0]     OE_DATA_64_const_net_13;
wire   [3:0]     OE_DATA_65_const_net_13;
wire   [3:0]     OE_DATA_66_const_net_13;
wire   [3:0]     OE_DATA_67_const_net_13;
wire   [3:0]     OE_DATA_68_const_net_13;
wire   [3:0]     OE_DATA_69_const_net_13;
wire   [3:0]     OE_DATA_70_const_net_13;
wire   [3:0]     OE_DATA_71_const_net_13;
wire   [3:0]     OE_DATA_72_const_net_13;
wire   [3:0]     OE_DATA_73_const_net_13;
wire   [3:0]     OE_DATA_74_const_net_13;
wire   [3:0]     OE_DATA_75_const_net_13;
wire   [3:0]     OE_DATA_76_const_net_13;
wire   [3:0]     OE_DATA_77_const_net_13;
wire   [3:0]     OE_DATA_78_const_net_13;
wire   [3:0]     OE_DATA_79_const_net_13;
wire   [3:0]     OE_DATA_80_const_net_13;
wire   [3:0]     OE_DATA_81_const_net_13;
wire   [3:0]     OE_DATA_82_const_net_13;
wire   [3:0]     OE_DATA_83_const_net_13;
wire   [3:0]     OE_DATA_84_const_net_13;
wire   [3:0]     OE_DATA_85_const_net_13;
wire   [3:0]     OE_DATA_86_const_net_13;
wire   [3:0]     OE_DATA_87_const_net_13;
wire   [3:0]     OE_DATA_88_const_net_13;
wire   [3:0]     OE_DATA_89_const_net_13;
wire   [3:0]     OE_DATA_90_const_net_13;
wire   [3:0]     OE_DATA_91_const_net_13;
wire   [3:0]     OE_DATA_92_const_net_13;
wire   [3:0]     OE_DATA_93_const_net_13;
wire   [3:0]     OE_DATA_94_const_net_13;
wire   [3:0]     OE_DATA_95_const_net_13;
wire   [3:0]     OE_DATA_96_const_net_13;
wire   [3:0]     OE_DATA_97_const_net_13;
wire   [3:0]     OE_DATA_98_const_net_13;
wire   [3:0]     OE_DATA_99_const_net_13;
wire   [3:0]     OE_DATA_100_const_net_13;
wire   [3:0]     OE_DATA_101_const_net_13;
wire   [3:0]     OE_DATA_102_const_net_13;
wire   [3:0]     OE_DATA_103_const_net_13;
wire   [3:0]     OE_DATA_104_const_net_13;
wire   [3:0]     OE_DATA_105_const_net_13;
wire   [3:0]     OE_DATA_106_const_net_13;
wire   [3:0]     OE_DATA_107_const_net_13;
wire   [3:0]     OE_DATA_108_const_net_13;
wire   [3:0]     OE_DATA_109_const_net_13;
wire   [3:0]     OE_DATA_110_const_net_13;
wire   [3:0]     OE_DATA_111_const_net_13;
wire   [3:0]     OE_DATA_112_const_net_13;
wire   [3:0]     OE_DATA_113_const_net_13;
wire   [3:0]     OE_DATA_114_const_net_13;
wire   [3:0]     OE_DATA_115_const_net_13;
wire   [3:0]     OE_DATA_116_const_net_13;
wire   [3:0]     OE_DATA_117_const_net_13;
wire   [3:0]     OE_DATA_118_const_net_13;
wire   [3:0]     OE_DATA_119_const_net_13;
wire   [3:0]     OE_DATA_120_const_net_13;
wire   [3:0]     OE_DATA_121_const_net_13;
wire   [3:0]     OE_DATA_122_const_net_13;
wire   [3:0]     OE_DATA_123_const_net_13;
wire   [3:0]     OE_DATA_124_const_net_13;
wire   [3:0]     OE_DATA_125_const_net_13;
wire   [3:0]     OE_DATA_126_const_net_13;
wire   [3:0]     OE_DATA_127_const_net_13;
wire   [1:0]     RX_DQS_90_const_net_14;
wire   [2:0]     FIFO_WR_PTR_const_net_14;
wire   [2:0]     FIFO_RD_PTR_const_net_14;
wire   [2:0]     EYE_MONITOR_LANE_WIDTH_const_net_14;
wire   [3:0]     TX_DATA_1_const_net_11;
wire   [3:0]     TX_DATA_2_const_net_13;
wire   [3:0]     TX_DATA_3_const_net_13;
wire   [3:0]     TX_DATA_4_const_net_13;
wire   [3:0]     TX_DATA_5_const_net_13;
wire   [3:0]     TX_DATA_6_const_net_13;
wire   [3:0]     TX_DATA_7_const_net_13;
wire   [3:0]     TX_DATA_8_const_net_13;
wire   [3:0]     TX_DATA_9_const_net_13;
wire   [3:0]     TX_DATA_10_const_net_13;
wire   [3:0]     TX_DATA_11_const_net_13;
wire   [3:0]     TX_DATA_12_const_net_14;
wire   [3:0]     TX_DATA_13_const_net_14;
wire   [3:0]     TX_DATA_14_const_net_14;
wire   [3:0]     TX_DATA_15_const_net_14;
wire   [3:0]     TX_DATA_16_const_net_14;
wire   [3:0]     TX_DATA_17_const_net_14;
wire   [3:0]     TX_DATA_18_const_net_14;
wire   [3:0]     TX_DATA_19_const_net_14;
wire   [3:0]     TX_DATA_20_const_net_14;
wire   [3:0]     TX_DATA_21_const_net_14;
wire   [3:0]     TX_DATA_22_const_net_14;
wire   [3:0]     TX_DATA_23_const_net_14;
wire   [3:0]     TX_DATA_24_const_net_14;
wire   [3:0]     TX_DATA_25_const_net_14;
wire   [3:0]     TX_DATA_26_const_net_14;
wire   [3:0]     TX_DATA_27_const_net_14;
wire   [3:0]     TX_DATA_28_const_net_14;
wire   [3:0]     TX_DATA_29_const_net_14;
wire   [3:0]     TX_DATA_30_const_net_14;
wire   [3:0]     TX_DATA_31_const_net_14;
wire   [3:0]     TX_DATA_32_const_net_14;
wire   [3:0]     TX_DATA_33_const_net_14;
wire   [3:0]     TX_DATA_34_const_net_14;
wire   [3:0]     TX_DATA_35_const_net_14;
wire   [3:0]     TX_DATA_36_const_net_14;
wire   [3:0]     TX_DATA_37_const_net_14;
wire   [3:0]     TX_DATA_38_const_net_14;
wire   [3:0]     TX_DATA_39_const_net_14;
wire   [3:0]     TX_DATA_40_const_net_14;
wire   [3:0]     TX_DATA_41_const_net_14;
wire   [3:0]     TX_DATA_42_const_net_14;
wire   [3:0]     TX_DATA_43_const_net_14;
wire   [3:0]     TX_DATA_44_const_net_14;
wire   [3:0]     TX_DATA_45_const_net_14;
wire   [3:0]     TX_DATA_46_const_net_14;
wire   [3:0]     TX_DATA_47_const_net_14;
wire   [3:0]     TX_DATA_48_const_net_14;
wire   [3:0]     TX_DATA_49_const_net_14;
wire   [3:0]     TX_DATA_50_const_net_14;
wire   [3:0]     TX_DATA_51_const_net_14;
wire   [3:0]     TX_DATA_52_const_net_14;
wire   [3:0]     TX_DATA_53_const_net_14;
wire   [3:0]     TX_DATA_54_const_net_14;
wire   [3:0]     TX_DATA_55_const_net_14;
wire   [3:0]     TX_DATA_56_const_net_14;
wire   [3:0]     TX_DATA_57_const_net_14;
wire   [3:0]     TX_DATA_58_const_net_14;
wire   [3:0]     TX_DATA_59_const_net_14;
wire   [3:0]     TX_DATA_60_const_net_14;
wire   [3:0]     TX_DATA_61_const_net_14;
wire   [3:0]     TX_DATA_62_const_net_14;
wire   [3:0]     TX_DATA_63_const_net_14;
wire   [3:0]     TX_DATA_64_const_net_14;
wire   [3:0]     TX_DATA_65_const_net_14;
wire   [3:0]     TX_DATA_66_const_net_14;
wire   [3:0]     TX_DATA_67_const_net_14;
wire   [3:0]     TX_DATA_68_const_net_14;
wire   [3:0]     TX_DATA_69_const_net_14;
wire   [3:0]     TX_DATA_70_const_net_14;
wire   [3:0]     TX_DATA_71_const_net_14;
wire   [3:0]     TX_DATA_72_const_net_14;
wire   [3:0]     TX_DATA_73_const_net_14;
wire   [3:0]     TX_DATA_74_const_net_14;
wire   [3:0]     TX_DATA_75_const_net_14;
wire   [3:0]     TX_DATA_76_const_net_14;
wire   [3:0]     TX_DATA_77_const_net_14;
wire   [3:0]     TX_DATA_78_const_net_14;
wire   [3:0]     TX_DATA_79_const_net_14;
wire   [3:0]     TX_DATA_80_const_net_14;
wire   [3:0]     TX_DATA_81_const_net_14;
wire   [3:0]     TX_DATA_82_const_net_14;
wire   [3:0]     TX_DATA_83_const_net_14;
wire   [3:0]     TX_DATA_84_const_net_14;
wire   [3:0]     TX_DATA_85_const_net_14;
wire   [3:0]     TX_DATA_86_const_net_14;
wire   [3:0]     TX_DATA_87_const_net_14;
wire   [3:0]     TX_DATA_88_const_net_14;
wire   [3:0]     TX_DATA_89_const_net_14;
wire   [3:0]     TX_DATA_90_const_net_14;
wire   [3:0]     TX_DATA_91_const_net_14;
wire   [3:0]     TX_DATA_92_const_net_14;
wire   [3:0]     TX_DATA_93_const_net_14;
wire   [3:0]     TX_DATA_94_const_net_14;
wire   [3:0]     TX_DATA_95_const_net_14;
wire   [3:0]     TX_DATA_96_const_net_14;
wire   [3:0]     TX_DATA_97_const_net_14;
wire   [3:0]     TX_DATA_98_const_net_14;
wire   [3:0]     TX_DATA_99_const_net_14;
wire   [3:0]     TX_DATA_100_const_net_14;
wire   [3:0]     TX_DATA_101_const_net_14;
wire   [3:0]     TX_DATA_102_const_net_14;
wire   [3:0]     TX_DATA_103_const_net_14;
wire   [3:0]     TX_DATA_104_const_net_14;
wire   [3:0]     TX_DATA_105_const_net_14;
wire   [3:0]     TX_DATA_106_const_net_14;
wire   [3:0]     TX_DATA_107_const_net_14;
wire   [3:0]     TX_DATA_108_const_net_14;
wire   [3:0]     TX_DATA_109_const_net_14;
wire   [3:0]     TX_DATA_110_const_net_14;
wire   [3:0]     TX_DATA_111_const_net_14;
wire   [3:0]     TX_DATA_112_const_net_14;
wire   [3:0]     TX_DATA_113_const_net_14;
wire   [3:0]     TX_DATA_114_const_net_14;
wire   [3:0]     TX_DATA_115_const_net_14;
wire   [3:0]     TX_DATA_116_const_net_14;
wire   [3:0]     TX_DATA_117_const_net_14;
wire   [3:0]     TX_DATA_118_const_net_14;
wire   [3:0]     TX_DATA_119_const_net_14;
wire   [3:0]     TX_DATA_120_const_net_14;
wire   [3:0]     TX_DATA_121_const_net_14;
wire   [3:0]     TX_DATA_122_const_net_14;
wire   [3:0]     TX_DATA_123_const_net_14;
wire   [3:0]     TX_DATA_124_const_net_14;
wire   [3:0]     TX_DATA_125_const_net_14;
wire   [3:0]     TX_DATA_126_const_net_14;
wire   [3:0]     TX_DATA_127_const_net_14;
wire   [3:0]     OE_DATA_1_const_net_14;
wire   [3:0]     OE_DATA_2_const_net_14;
wire   [3:0]     OE_DATA_3_const_net_14;
wire   [3:0]     OE_DATA_4_const_net_14;
wire   [3:0]     OE_DATA_5_const_net_14;
wire   [3:0]     OE_DATA_6_const_net_14;
wire   [3:0]     OE_DATA_7_const_net_14;
wire   [3:0]     OE_DATA_8_const_net_14;
wire   [3:0]     OE_DATA_9_const_net_14;
wire   [3:0]     OE_DATA_10_const_net_14;
wire   [3:0]     OE_DATA_11_const_net_14;
wire   [3:0]     OE_DATA_12_const_net_14;
wire   [3:0]     OE_DATA_13_const_net_14;
wire   [3:0]     OE_DATA_14_const_net_14;
wire   [3:0]     OE_DATA_15_const_net_14;
wire   [3:0]     OE_DATA_16_const_net_14;
wire   [3:0]     OE_DATA_17_const_net_14;
wire   [3:0]     OE_DATA_18_const_net_14;
wire   [3:0]     OE_DATA_19_const_net_14;
wire   [3:0]     OE_DATA_20_const_net_14;
wire   [3:0]     OE_DATA_21_const_net_14;
wire   [3:0]     OE_DATA_22_const_net_14;
wire   [3:0]     OE_DATA_23_const_net_14;
wire   [3:0]     OE_DATA_24_const_net_14;
wire   [3:0]     OE_DATA_25_const_net_14;
wire   [3:0]     OE_DATA_26_const_net_14;
wire   [3:0]     OE_DATA_27_const_net_14;
wire   [3:0]     OE_DATA_28_const_net_14;
wire   [3:0]     OE_DATA_29_const_net_14;
wire   [3:0]     OE_DATA_30_const_net_14;
wire   [3:0]     OE_DATA_31_const_net_14;
wire   [3:0]     OE_DATA_32_const_net_14;
wire   [3:0]     OE_DATA_33_const_net_14;
wire   [3:0]     OE_DATA_34_const_net_14;
wire   [3:0]     OE_DATA_35_const_net_14;
wire   [3:0]     OE_DATA_36_const_net_14;
wire   [3:0]     OE_DATA_37_const_net_14;
wire   [3:0]     OE_DATA_38_const_net_14;
wire   [3:0]     OE_DATA_39_const_net_14;
wire   [3:0]     OE_DATA_40_const_net_14;
wire   [3:0]     OE_DATA_41_const_net_14;
wire   [3:0]     OE_DATA_42_const_net_14;
wire   [3:0]     OE_DATA_43_const_net_14;
wire   [3:0]     OE_DATA_44_const_net_14;
wire   [3:0]     OE_DATA_45_const_net_14;
wire   [3:0]     OE_DATA_46_const_net_14;
wire   [3:0]     OE_DATA_47_const_net_14;
wire   [3:0]     OE_DATA_48_const_net_14;
wire   [3:0]     OE_DATA_49_const_net_14;
wire   [3:0]     OE_DATA_50_const_net_14;
wire   [3:0]     OE_DATA_51_const_net_14;
wire   [3:0]     OE_DATA_52_const_net_14;
wire   [3:0]     OE_DATA_53_const_net_14;
wire   [3:0]     OE_DATA_54_const_net_14;
wire   [3:0]     OE_DATA_55_const_net_14;
wire   [3:0]     OE_DATA_56_const_net_14;
wire   [3:0]     OE_DATA_57_const_net_14;
wire   [3:0]     OE_DATA_58_const_net_14;
wire   [3:0]     OE_DATA_59_const_net_14;
wire   [3:0]     OE_DATA_60_const_net_14;
wire   [3:0]     OE_DATA_61_const_net_14;
wire   [3:0]     OE_DATA_62_const_net_14;
wire   [3:0]     OE_DATA_63_const_net_14;
wire   [3:0]     OE_DATA_64_const_net_14;
wire   [3:0]     OE_DATA_65_const_net_14;
wire   [3:0]     OE_DATA_66_const_net_14;
wire   [3:0]     OE_DATA_67_const_net_14;
wire   [3:0]     OE_DATA_68_const_net_14;
wire   [3:0]     OE_DATA_69_const_net_14;
wire   [3:0]     OE_DATA_70_const_net_14;
wire   [3:0]     OE_DATA_71_const_net_14;
wire   [3:0]     OE_DATA_72_const_net_14;
wire   [3:0]     OE_DATA_73_const_net_14;
wire   [3:0]     OE_DATA_74_const_net_14;
wire   [3:0]     OE_DATA_75_const_net_14;
wire   [3:0]     OE_DATA_76_const_net_14;
wire   [3:0]     OE_DATA_77_const_net_14;
wire   [3:0]     OE_DATA_78_const_net_14;
wire   [3:0]     OE_DATA_79_const_net_14;
wire   [3:0]     OE_DATA_80_const_net_14;
wire   [3:0]     OE_DATA_81_const_net_14;
wire   [3:0]     OE_DATA_82_const_net_14;
wire   [3:0]     OE_DATA_83_const_net_14;
wire   [3:0]     OE_DATA_84_const_net_14;
wire   [3:0]     OE_DATA_85_const_net_14;
wire   [3:0]     OE_DATA_86_const_net_14;
wire   [3:0]     OE_DATA_87_const_net_14;
wire   [3:0]     OE_DATA_88_const_net_14;
wire   [3:0]     OE_DATA_89_const_net_14;
wire   [3:0]     OE_DATA_90_const_net_14;
wire   [3:0]     OE_DATA_91_const_net_14;
wire   [3:0]     OE_DATA_92_const_net_14;
wire   [3:0]     OE_DATA_93_const_net_14;
wire   [3:0]     OE_DATA_94_const_net_14;
wire   [3:0]     OE_DATA_95_const_net_14;
wire   [3:0]     OE_DATA_96_const_net_14;
wire   [3:0]     OE_DATA_97_const_net_14;
wire   [3:0]     OE_DATA_98_const_net_14;
wire   [3:0]     OE_DATA_99_const_net_14;
wire   [3:0]     OE_DATA_100_const_net_14;
wire   [3:0]     OE_DATA_101_const_net_14;
wire   [3:0]     OE_DATA_102_const_net_14;
wire   [3:0]     OE_DATA_103_const_net_14;
wire   [3:0]     OE_DATA_104_const_net_14;
wire   [3:0]     OE_DATA_105_const_net_14;
wire   [3:0]     OE_DATA_106_const_net_14;
wire   [3:0]     OE_DATA_107_const_net_14;
wire   [3:0]     OE_DATA_108_const_net_14;
wire   [3:0]     OE_DATA_109_const_net_14;
wire   [3:0]     OE_DATA_110_const_net_14;
wire   [3:0]     OE_DATA_111_const_net_14;
wire   [3:0]     OE_DATA_112_const_net_14;
wire   [3:0]     OE_DATA_113_const_net_14;
wire   [3:0]     OE_DATA_114_const_net_14;
wire   [3:0]     OE_DATA_115_const_net_14;
wire   [3:0]     OE_DATA_116_const_net_14;
wire   [3:0]     OE_DATA_117_const_net_14;
wire   [3:0]     OE_DATA_118_const_net_14;
wire   [3:0]     OE_DATA_119_const_net_14;
wire   [3:0]     OE_DATA_120_const_net_14;
wire   [3:0]     OE_DATA_121_const_net_14;
wire   [3:0]     OE_DATA_122_const_net_14;
wire   [3:0]     OE_DATA_123_const_net_14;
wire   [3:0]     OE_DATA_124_const_net_14;
wire   [3:0]     OE_DATA_125_const_net_14;
wire   [3:0]     OE_DATA_126_const_net_14;
wire   [3:0]     OE_DATA_127_const_net_14;
wire   [10:0]    CDR_CLK_B_SEL_const_net_0;
wire   [2:0]     FIFO_WR_PTR_const_net_15;
wire   [2:0]     FIFO_RD_PTR_const_net_15;
wire   [2:0]     EYE_MONITOR_LANE_WIDTH_const_net_15;
wire   [7:0]     TX_DATA_1_const_net_12;
wire   [7:0]     TX_DATA_2_const_net_14;
wire   [7:0]     TX_DATA_3_const_net_14;
wire   [7:0]     TX_DATA_4_const_net_14;
wire   [7:0]     TX_DATA_5_const_net_14;
wire   [7:0]     TX_DATA_6_const_net_14;
wire   [7:0]     TX_DATA_7_const_net_14;
wire   [7:0]     TX_DATA_8_const_net_14;
wire   [7:0]     TX_DATA_9_const_net_14;
wire   [7:0]     TX_DATA_10_const_net_14;
wire   [7:0]     TX_DATA_11_const_net_14;
wire   [7:0]     TX_DATA_12_const_net_15;
wire   [7:0]     TX_DATA_13_const_net_15;
wire   [7:0]     TX_DATA_14_const_net_15;
wire   [7:0]     TX_DATA_15_const_net_15;
wire   [7:0]     TX_DATA_16_const_net_15;
wire   [7:0]     TX_DATA_17_const_net_15;
wire   [7:0]     TX_DATA_18_const_net_15;
wire   [7:0]     TX_DATA_19_const_net_15;
wire   [7:0]     TX_DATA_20_const_net_15;
wire   [7:0]     TX_DATA_21_const_net_15;
wire   [7:0]     TX_DATA_22_const_net_15;
wire   [7:0]     TX_DATA_23_const_net_15;
wire   [7:0]     TX_DATA_24_const_net_15;
wire   [7:0]     TX_DATA_25_const_net_15;
wire   [7:0]     TX_DATA_26_const_net_15;
wire   [7:0]     TX_DATA_27_const_net_15;
wire   [7:0]     TX_DATA_28_const_net_15;
wire   [7:0]     TX_DATA_29_const_net_15;
wire   [7:0]     TX_DATA_30_const_net_15;
wire   [7:0]     TX_DATA_31_const_net_15;
wire   [7:0]     TX_DATA_32_const_net_15;
wire   [7:0]     TX_DATA_33_const_net_15;
wire   [7:0]     TX_DATA_34_const_net_15;
wire   [7:0]     TX_DATA_35_const_net_15;
wire   [7:0]     TX_DATA_36_const_net_15;
wire   [7:0]     TX_DATA_37_const_net_15;
wire   [7:0]     TX_DATA_38_const_net_15;
wire   [7:0]     TX_DATA_39_const_net_15;
wire   [7:0]     TX_DATA_40_const_net_15;
wire   [7:0]     TX_DATA_41_const_net_15;
wire   [7:0]     TX_DATA_42_const_net_15;
wire   [7:0]     TX_DATA_43_const_net_15;
wire   [7:0]     TX_DATA_44_const_net_15;
wire   [7:0]     TX_DATA_45_const_net_15;
wire   [7:0]     TX_DATA_46_const_net_15;
wire   [7:0]     TX_DATA_47_const_net_15;
wire   [7:0]     TX_DATA_48_const_net_15;
wire   [7:0]     TX_DATA_49_const_net_15;
wire   [7:0]     TX_DATA_50_const_net_15;
wire   [7:0]     TX_DATA_51_const_net_15;
wire   [7:0]     TX_DATA_52_const_net_15;
wire   [7:0]     TX_DATA_53_const_net_15;
wire   [7:0]     TX_DATA_54_const_net_15;
wire   [7:0]     TX_DATA_55_const_net_15;
wire   [7:0]     TX_DATA_56_const_net_15;
wire   [7:0]     TX_DATA_57_const_net_15;
wire   [7:0]     TX_DATA_58_const_net_15;
wire   [7:0]     TX_DATA_59_const_net_15;
wire   [7:0]     TX_DATA_60_const_net_15;
wire   [7:0]     TX_DATA_61_const_net_15;
wire   [7:0]     TX_DATA_62_const_net_15;
wire   [7:0]     TX_DATA_63_const_net_15;
wire   [7:0]     TX_DATA_64_const_net_15;
wire   [7:0]     TX_DATA_65_const_net_15;
wire   [7:0]     TX_DATA_66_const_net_15;
wire   [7:0]     TX_DATA_67_const_net_15;
wire   [7:0]     TX_DATA_68_const_net_15;
wire   [7:0]     TX_DATA_69_const_net_15;
wire   [7:0]     TX_DATA_70_const_net_15;
wire   [7:0]     TX_DATA_71_const_net_15;
wire   [7:0]     TX_DATA_72_const_net_15;
wire   [7:0]     TX_DATA_73_const_net_15;
wire   [7:0]     TX_DATA_74_const_net_15;
wire   [7:0]     TX_DATA_75_const_net_15;
wire   [7:0]     TX_DATA_76_const_net_15;
wire   [7:0]     TX_DATA_77_const_net_15;
wire   [7:0]     TX_DATA_78_const_net_15;
wire   [7:0]     TX_DATA_79_const_net_15;
wire   [7:0]     TX_DATA_80_const_net_15;
wire   [7:0]     TX_DATA_81_const_net_15;
wire   [7:0]     TX_DATA_82_const_net_15;
wire   [7:0]     TX_DATA_83_const_net_15;
wire   [7:0]     TX_DATA_84_const_net_15;
wire   [7:0]     TX_DATA_85_const_net_15;
wire   [7:0]     TX_DATA_86_const_net_15;
wire   [7:0]     TX_DATA_87_const_net_15;
wire   [7:0]     TX_DATA_88_const_net_15;
wire   [7:0]     TX_DATA_89_const_net_15;
wire   [7:0]     TX_DATA_90_const_net_15;
wire   [7:0]     TX_DATA_91_const_net_15;
wire   [7:0]     TX_DATA_92_const_net_15;
wire   [7:0]     TX_DATA_93_const_net_15;
wire   [7:0]     TX_DATA_94_const_net_15;
wire   [7:0]     TX_DATA_95_const_net_15;
wire   [7:0]     TX_DATA_96_const_net_15;
wire   [7:0]     TX_DATA_97_const_net_15;
wire   [7:0]     TX_DATA_98_const_net_15;
wire   [7:0]     TX_DATA_99_const_net_15;
wire   [7:0]     TX_DATA_100_const_net_15;
wire   [7:0]     TX_DATA_101_const_net_15;
wire   [7:0]     TX_DATA_102_const_net_15;
wire   [7:0]     TX_DATA_103_const_net_15;
wire   [7:0]     TX_DATA_104_const_net_15;
wire   [7:0]     TX_DATA_105_const_net_15;
wire   [7:0]     TX_DATA_106_const_net_15;
wire   [7:0]     TX_DATA_107_const_net_15;
wire   [7:0]     TX_DATA_108_const_net_15;
wire   [7:0]     TX_DATA_109_const_net_15;
wire   [7:0]     TX_DATA_110_const_net_15;
wire   [7:0]     TX_DATA_111_const_net_15;
wire   [7:0]     TX_DATA_112_const_net_15;
wire   [7:0]     TX_DATA_113_const_net_15;
wire   [7:0]     TX_DATA_114_const_net_15;
wire   [7:0]     TX_DATA_115_const_net_15;
wire   [7:0]     TX_DATA_116_const_net_15;
wire   [7:0]     TX_DATA_117_const_net_15;
wire   [7:0]     TX_DATA_118_const_net_15;
wire   [7:0]     TX_DATA_119_const_net_15;
wire   [7:0]     TX_DATA_120_const_net_15;
wire   [7:0]     TX_DATA_121_const_net_15;
wire   [7:0]     TX_DATA_122_const_net_15;
wire   [7:0]     TX_DATA_123_const_net_15;
wire   [7:0]     TX_DATA_124_const_net_15;
wire   [7:0]     TX_DATA_125_const_net_15;
wire   [7:0]     TX_DATA_126_const_net_15;
wire   [7:0]     TX_DATA_127_const_net_15;
wire   [3:0]     OE_DATA_1_const_net_15;
wire   [3:0]     OE_DATA_2_const_net_15;
wire   [3:0]     OE_DATA_3_const_net_15;
wire   [3:0]     OE_DATA_4_const_net_15;
wire   [3:0]     OE_DATA_5_const_net_15;
wire   [3:0]     OE_DATA_6_const_net_15;
wire   [3:0]     OE_DATA_7_const_net_15;
wire   [3:0]     OE_DATA_8_const_net_15;
wire   [3:0]     OE_DATA_9_const_net_15;
wire   [3:0]     OE_DATA_10_const_net_15;
wire   [3:0]     OE_DATA_11_const_net_15;
wire   [3:0]     OE_DATA_12_const_net_15;
wire   [3:0]     OE_DATA_13_const_net_15;
wire   [3:0]     OE_DATA_14_const_net_15;
wire   [3:0]     OE_DATA_15_const_net_15;
wire   [3:0]     OE_DATA_16_const_net_15;
wire   [3:0]     OE_DATA_17_const_net_15;
wire   [3:0]     OE_DATA_18_const_net_15;
wire   [3:0]     OE_DATA_19_const_net_15;
wire   [3:0]     OE_DATA_20_const_net_15;
wire   [3:0]     OE_DATA_21_const_net_15;
wire   [3:0]     OE_DATA_22_const_net_15;
wire   [3:0]     OE_DATA_23_const_net_15;
wire   [3:0]     OE_DATA_24_const_net_15;
wire   [3:0]     OE_DATA_25_const_net_15;
wire   [3:0]     OE_DATA_26_const_net_15;
wire   [3:0]     OE_DATA_27_const_net_15;
wire   [3:0]     OE_DATA_28_const_net_15;
wire   [3:0]     OE_DATA_29_const_net_15;
wire   [3:0]     OE_DATA_30_const_net_15;
wire   [3:0]     OE_DATA_31_const_net_15;
wire   [3:0]     OE_DATA_32_const_net_15;
wire   [3:0]     OE_DATA_33_const_net_15;
wire   [3:0]     OE_DATA_34_const_net_15;
wire   [3:0]     OE_DATA_35_const_net_15;
wire   [3:0]     OE_DATA_36_const_net_15;
wire   [3:0]     OE_DATA_37_const_net_15;
wire   [3:0]     OE_DATA_38_const_net_15;
wire   [3:0]     OE_DATA_39_const_net_15;
wire   [3:0]     OE_DATA_40_const_net_15;
wire   [3:0]     OE_DATA_41_const_net_15;
wire   [3:0]     OE_DATA_42_const_net_15;
wire   [3:0]     OE_DATA_43_const_net_15;
wire   [3:0]     OE_DATA_44_const_net_15;
wire   [3:0]     OE_DATA_45_const_net_15;
wire   [3:0]     OE_DATA_46_const_net_15;
wire   [3:0]     OE_DATA_47_const_net_15;
wire   [3:0]     OE_DATA_48_const_net_15;
wire   [3:0]     OE_DATA_49_const_net_15;
wire   [3:0]     OE_DATA_50_const_net_15;
wire   [3:0]     OE_DATA_51_const_net_15;
wire   [3:0]     OE_DATA_52_const_net_15;
wire   [3:0]     OE_DATA_53_const_net_15;
wire   [3:0]     OE_DATA_54_const_net_15;
wire   [3:0]     OE_DATA_55_const_net_15;
wire   [3:0]     OE_DATA_56_const_net_15;
wire   [3:0]     OE_DATA_57_const_net_15;
wire   [3:0]     OE_DATA_58_const_net_15;
wire   [3:0]     OE_DATA_59_const_net_15;
wire   [3:0]     OE_DATA_60_const_net_15;
wire   [3:0]     OE_DATA_61_const_net_15;
wire   [3:0]     OE_DATA_62_const_net_15;
wire   [3:0]     OE_DATA_63_const_net_15;
wire   [3:0]     OE_DATA_64_const_net_15;
wire   [3:0]     OE_DATA_65_const_net_15;
wire   [3:0]     OE_DATA_66_const_net_15;
wire   [3:0]     OE_DATA_67_const_net_15;
wire   [3:0]     OE_DATA_68_const_net_15;
wire   [3:0]     OE_DATA_69_const_net_15;
wire   [3:0]     OE_DATA_70_const_net_15;
wire   [3:0]     OE_DATA_71_const_net_15;
wire   [3:0]     OE_DATA_72_const_net_15;
wire   [3:0]     OE_DATA_73_const_net_15;
wire   [3:0]     OE_DATA_74_const_net_15;
wire   [3:0]     OE_DATA_75_const_net_15;
wire   [3:0]     OE_DATA_76_const_net_15;
wire   [3:0]     OE_DATA_77_const_net_15;
wire   [3:0]     OE_DATA_78_const_net_15;
wire   [3:0]     OE_DATA_79_const_net_15;
wire   [3:0]     OE_DATA_80_const_net_15;
wire   [3:0]     OE_DATA_81_const_net_15;
wire   [3:0]     OE_DATA_82_const_net_15;
wire   [3:0]     OE_DATA_83_const_net_15;
wire   [3:0]     OE_DATA_84_const_net_15;
wire   [3:0]     OE_DATA_85_const_net_15;
wire   [3:0]     OE_DATA_86_const_net_15;
wire   [3:0]     OE_DATA_87_const_net_15;
wire   [3:0]     OE_DATA_88_const_net_15;
wire   [3:0]     OE_DATA_89_const_net_15;
wire   [3:0]     OE_DATA_90_const_net_15;
wire   [3:0]     OE_DATA_91_const_net_15;
wire   [3:0]     OE_DATA_92_const_net_15;
wire   [3:0]     OE_DATA_93_const_net_15;
wire   [3:0]     OE_DATA_94_const_net_15;
wire   [3:0]     OE_DATA_95_const_net_15;
wire   [3:0]     OE_DATA_96_const_net_15;
wire   [3:0]     OE_DATA_97_const_net_15;
wire   [3:0]     OE_DATA_98_const_net_15;
wire   [3:0]     OE_DATA_99_const_net_15;
wire   [3:0]     OE_DATA_100_const_net_15;
wire   [3:0]     OE_DATA_101_const_net_15;
wire   [3:0]     OE_DATA_102_const_net_15;
wire   [3:0]     OE_DATA_103_const_net_15;
wire   [3:0]     OE_DATA_104_const_net_15;
wire   [3:0]     OE_DATA_105_const_net_15;
wire   [3:0]     OE_DATA_106_const_net_15;
wire   [3:0]     OE_DATA_107_const_net_15;
wire   [3:0]     OE_DATA_108_const_net_15;
wire   [3:0]     OE_DATA_109_const_net_15;
wire   [3:0]     OE_DATA_110_const_net_15;
wire   [3:0]     OE_DATA_111_const_net_15;
wire   [3:0]     OE_DATA_112_const_net_15;
wire   [3:0]     OE_DATA_113_const_net_15;
wire   [3:0]     OE_DATA_114_const_net_15;
wire   [3:0]     OE_DATA_115_const_net_15;
wire   [3:0]     OE_DATA_116_const_net_15;
wire   [3:0]     OE_DATA_117_const_net_15;
wire   [3:0]     OE_DATA_118_const_net_15;
wire   [3:0]     OE_DATA_119_const_net_15;
wire   [3:0]     OE_DATA_120_const_net_15;
wire   [3:0]     OE_DATA_121_const_net_15;
wire   [3:0]     OE_DATA_122_const_net_15;
wire   [3:0]     OE_DATA_123_const_net_15;
wire   [3:0]     OE_DATA_124_const_net_15;
wire   [3:0]     OE_DATA_125_const_net_15;
wire   [3:0]     OE_DATA_126_const_net_15;
wire   [3:0]     OE_DATA_127_const_net_15;
wire   [7:0]     TX_DATA_8_const_net_15;
wire   [7:0]     TX_DATA_9_const_net_15;
wire   [7:0]     TX_DATA_10_const_net_15;
wire   [7:0]     TX_DATA_11_const_net_15;
wire   [7:0]     TX_DATA_12_const_net_16;
wire   [7:0]     TX_DATA_13_const_net_16;
wire   [7:0]     TX_DATA_14_const_net_16;
wire   [7:0]     TX_DATA_15_const_net_16;
wire   [7:0]     TX_DATA_16_const_net_16;
wire   [7:0]     TX_DATA_17_const_net_16;
wire   [7:0]     TX_DATA_18_const_net_16;
wire   [7:0]     TX_DATA_19_const_net_16;
wire   [7:0]     TX_DATA_20_const_net_16;
wire   [7:0]     TX_DATA_21_const_net_16;
wire   [7:0]     TX_DATA_22_const_net_16;
wire   [7:0]     TX_DATA_23_const_net_16;
wire   [7:0]     TX_DATA_24_const_net_16;
wire   [7:0]     TX_DATA_25_const_net_16;
wire   [7:0]     TX_DATA_26_const_net_16;
wire   [7:0]     TX_DATA_27_const_net_16;
wire   [7:0]     TX_DATA_28_const_net_16;
wire   [7:0]     TX_DATA_29_const_net_16;
wire   [7:0]     TX_DATA_30_const_net_16;
wire   [7:0]     TX_DATA_31_const_net_16;
wire   [7:0]     TX_DATA_32_const_net_16;
wire   [7:0]     TX_DATA_33_const_net_16;
wire   [7:0]     TX_DATA_34_const_net_16;
wire   [7:0]     TX_DATA_35_const_net_16;
wire   [7:0]     TX_DATA_36_const_net_16;
wire   [7:0]     TX_DATA_37_const_net_16;
wire   [7:0]     TX_DATA_38_const_net_16;
wire   [7:0]     TX_DATA_39_const_net_16;
wire   [7:0]     TX_DATA_40_const_net_16;
wire   [7:0]     TX_DATA_41_const_net_16;
wire   [7:0]     TX_DATA_42_const_net_16;
wire   [7:0]     TX_DATA_43_const_net_16;
wire   [7:0]     TX_DATA_44_const_net_16;
wire   [7:0]     TX_DATA_45_const_net_16;
wire   [7:0]     TX_DATA_46_const_net_16;
wire   [7:0]     TX_DATA_47_const_net_16;
wire   [7:0]     TX_DATA_48_const_net_16;
wire   [7:0]     TX_DATA_49_const_net_16;
wire   [7:0]     TX_DATA_50_const_net_16;
wire   [7:0]     TX_DATA_51_const_net_16;
wire   [7:0]     TX_DATA_52_const_net_16;
wire   [7:0]     TX_DATA_53_const_net_16;
wire   [7:0]     TX_DATA_54_const_net_16;
wire   [7:0]     TX_DATA_55_const_net_16;
wire   [7:0]     TX_DATA_56_const_net_16;
wire   [7:0]     TX_DATA_57_const_net_16;
wire   [7:0]     TX_DATA_58_const_net_16;
wire   [7:0]     TX_DATA_59_const_net_16;
wire   [7:0]     TX_DATA_60_const_net_16;
wire   [7:0]     TX_DATA_61_const_net_16;
wire   [7:0]     TX_DATA_62_const_net_16;
wire   [7:0]     TX_DATA_63_const_net_16;
wire   [7:0]     TX_DATA_64_const_net_16;
wire   [7:0]     TX_DATA_65_const_net_16;
wire   [7:0]     TX_DATA_66_const_net_16;
wire   [7:0]     TX_DATA_67_const_net_16;
wire   [7:0]     TX_DATA_68_const_net_16;
wire   [7:0]     TX_DATA_69_const_net_16;
wire   [7:0]     TX_DATA_70_const_net_16;
wire   [7:0]     TX_DATA_71_const_net_16;
wire   [7:0]     TX_DATA_72_const_net_16;
wire   [7:0]     TX_DATA_73_const_net_16;
wire   [7:0]     TX_DATA_74_const_net_16;
wire   [7:0]     TX_DATA_75_const_net_16;
wire   [7:0]     TX_DATA_76_const_net_16;
wire   [7:0]     TX_DATA_77_const_net_16;
wire   [7:0]     TX_DATA_78_const_net_16;
wire   [7:0]     TX_DATA_79_const_net_16;
wire   [7:0]     TX_DATA_80_const_net_16;
wire   [7:0]     TX_DATA_81_const_net_16;
wire   [7:0]     TX_DATA_82_const_net_16;
wire   [7:0]     TX_DATA_83_const_net_16;
wire   [7:0]     TX_DATA_84_const_net_16;
wire   [7:0]     TX_DATA_85_const_net_16;
wire   [7:0]     TX_DATA_86_const_net_16;
wire   [7:0]     TX_DATA_87_const_net_16;
wire   [7:0]     TX_DATA_88_const_net_16;
wire   [7:0]     TX_DATA_89_const_net_16;
wire   [7:0]     TX_DATA_90_const_net_16;
wire   [7:0]     TX_DATA_91_const_net_16;
wire   [7:0]     TX_DATA_92_const_net_16;
wire   [7:0]     TX_DATA_93_const_net_16;
wire   [7:0]     TX_DATA_94_const_net_16;
wire   [7:0]     TX_DATA_95_const_net_16;
wire   [7:0]     TX_DATA_96_const_net_16;
wire   [7:0]     TX_DATA_97_const_net_16;
wire   [7:0]     TX_DATA_98_const_net_16;
wire   [7:0]     TX_DATA_99_const_net_16;
wire   [7:0]     TX_DATA_100_const_net_16;
wire   [7:0]     TX_DATA_101_const_net_16;
wire   [7:0]     TX_DATA_102_const_net_16;
wire   [7:0]     TX_DATA_103_const_net_16;
wire   [7:0]     TX_DATA_104_const_net_16;
wire   [7:0]     TX_DATA_105_const_net_16;
wire   [7:0]     TX_DATA_106_const_net_16;
wire   [7:0]     TX_DATA_107_const_net_16;
wire   [7:0]     TX_DATA_108_const_net_16;
wire   [7:0]     TX_DATA_109_const_net_16;
wire   [7:0]     TX_DATA_110_const_net_16;
wire   [7:0]     TX_DATA_111_const_net_16;
wire   [7:0]     TX_DATA_112_const_net_16;
wire   [7:0]     TX_DATA_113_const_net_16;
wire   [7:0]     TX_DATA_114_const_net_16;
wire   [7:0]     TX_DATA_115_const_net_16;
wire   [7:0]     TX_DATA_116_const_net_16;
wire   [7:0]     TX_DATA_117_const_net_16;
wire   [7:0]     TX_DATA_118_const_net_16;
wire   [7:0]     TX_DATA_119_const_net_16;
wire   [7:0]     TX_DATA_120_const_net_16;
wire   [7:0]     TX_DATA_121_const_net_16;
wire   [7:0]     TX_DATA_122_const_net_16;
wire   [7:0]     TX_DATA_123_const_net_16;
wire   [7:0]     TX_DATA_124_const_net_16;
wire   [7:0]     TX_DATA_125_const_net_16;
wire   [7:0]     TX_DATA_126_const_net_16;
wire   [7:0]     TX_DATA_127_const_net_16;
wire   [3:0]     OE_DATA_8_const_net_16;
wire   [3:0]     OE_DATA_9_const_net_16;
wire   [3:0]     OE_DATA_10_const_net_16;
wire   [3:0]     OE_DATA_11_const_net_16;
wire   [3:0]     OE_DATA_12_const_net_16;
wire   [3:0]     OE_DATA_13_const_net_16;
wire   [3:0]     OE_DATA_14_const_net_16;
wire   [3:0]     OE_DATA_15_const_net_16;
wire   [3:0]     OE_DATA_16_const_net_16;
wire   [3:0]     OE_DATA_17_const_net_16;
wire   [3:0]     OE_DATA_18_const_net_16;
wire   [3:0]     OE_DATA_19_const_net_16;
wire   [3:0]     OE_DATA_20_const_net_16;
wire   [3:0]     OE_DATA_21_const_net_16;
wire   [3:0]     OE_DATA_22_const_net_16;
wire   [3:0]     OE_DATA_23_const_net_16;
wire   [3:0]     OE_DATA_24_const_net_16;
wire   [3:0]     OE_DATA_25_const_net_16;
wire   [3:0]     OE_DATA_26_const_net_16;
wire   [3:0]     OE_DATA_27_const_net_16;
wire   [3:0]     OE_DATA_28_const_net_16;
wire   [3:0]     OE_DATA_29_const_net_16;
wire   [3:0]     OE_DATA_30_const_net_16;
wire   [3:0]     OE_DATA_31_const_net_16;
wire   [3:0]     OE_DATA_32_const_net_16;
wire   [3:0]     OE_DATA_33_const_net_16;
wire   [3:0]     OE_DATA_34_const_net_16;
wire   [3:0]     OE_DATA_35_const_net_16;
wire   [3:0]     OE_DATA_36_const_net_16;
wire   [3:0]     OE_DATA_37_const_net_16;
wire   [3:0]     OE_DATA_38_const_net_16;
wire   [3:0]     OE_DATA_39_const_net_16;
wire   [3:0]     OE_DATA_40_const_net_16;
wire   [3:0]     OE_DATA_41_const_net_16;
wire   [3:0]     OE_DATA_42_const_net_16;
wire   [3:0]     OE_DATA_43_const_net_16;
wire   [3:0]     OE_DATA_44_const_net_16;
wire   [3:0]     OE_DATA_45_const_net_16;
wire   [3:0]     OE_DATA_46_const_net_16;
wire   [3:0]     OE_DATA_47_const_net_16;
wire   [3:0]     OE_DATA_48_const_net_16;
wire   [3:0]     OE_DATA_49_const_net_16;
wire   [3:0]     OE_DATA_50_const_net_16;
wire   [3:0]     OE_DATA_51_const_net_16;
wire   [3:0]     OE_DATA_52_const_net_16;
wire   [3:0]     OE_DATA_53_const_net_16;
wire   [3:0]     OE_DATA_54_const_net_16;
wire   [3:0]     OE_DATA_55_const_net_16;
wire   [3:0]     OE_DATA_56_const_net_16;
wire   [3:0]     OE_DATA_57_const_net_16;
wire   [3:0]     OE_DATA_58_const_net_16;
wire   [3:0]     OE_DATA_59_const_net_16;
wire   [3:0]     OE_DATA_60_const_net_16;
wire   [3:0]     OE_DATA_61_const_net_16;
wire   [3:0]     OE_DATA_62_const_net_16;
wire   [3:0]     OE_DATA_63_const_net_16;
wire   [3:0]     OE_DATA_64_const_net_16;
wire   [3:0]     OE_DATA_65_const_net_16;
wire   [3:0]     OE_DATA_66_const_net_16;
wire   [3:0]     OE_DATA_67_const_net_16;
wire   [3:0]     OE_DATA_68_const_net_16;
wire   [3:0]     OE_DATA_69_const_net_16;
wire   [3:0]     OE_DATA_70_const_net_16;
wire   [3:0]     OE_DATA_71_const_net_16;
wire   [3:0]     OE_DATA_72_const_net_16;
wire   [3:0]     OE_DATA_73_const_net_16;
wire   [3:0]     OE_DATA_74_const_net_16;
wire   [3:0]     OE_DATA_75_const_net_16;
wire   [3:0]     OE_DATA_76_const_net_16;
wire   [3:0]     OE_DATA_77_const_net_16;
wire   [3:0]     OE_DATA_78_const_net_16;
wire   [3:0]     OE_DATA_79_const_net_16;
wire   [3:0]     OE_DATA_80_const_net_16;
wire   [3:0]     OE_DATA_81_const_net_16;
wire   [3:0]     OE_DATA_82_const_net_16;
wire   [3:0]     OE_DATA_83_const_net_16;
wire   [3:0]     OE_DATA_84_const_net_16;
wire   [3:0]     OE_DATA_85_const_net_16;
wire   [3:0]     OE_DATA_86_const_net_16;
wire   [3:0]     OE_DATA_87_const_net_16;
wire   [3:0]     OE_DATA_88_const_net_16;
wire   [3:0]     OE_DATA_89_const_net_16;
wire   [3:0]     OE_DATA_90_const_net_16;
wire   [3:0]     OE_DATA_91_const_net_16;
wire   [3:0]     OE_DATA_92_const_net_16;
wire   [3:0]     OE_DATA_93_const_net_16;
wire   [3:0]     OE_DATA_94_const_net_16;
wire   [3:0]     OE_DATA_95_const_net_16;
wire   [3:0]     OE_DATA_96_const_net_16;
wire   [3:0]     OE_DATA_97_const_net_16;
wire   [3:0]     OE_DATA_98_const_net_16;
wire   [3:0]     OE_DATA_99_const_net_16;
wire   [3:0]     OE_DATA_100_const_net_16;
wire   [3:0]     OE_DATA_101_const_net_16;
wire   [3:0]     OE_DATA_102_const_net_16;
wire   [3:0]     OE_DATA_103_const_net_16;
wire   [3:0]     OE_DATA_104_const_net_16;
wire   [3:0]     OE_DATA_105_const_net_16;
wire   [3:0]     OE_DATA_106_const_net_16;
wire   [3:0]     OE_DATA_107_const_net_16;
wire   [3:0]     OE_DATA_108_const_net_16;
wire   [3:0]     OE_DATA_109_const_net_16;
wire   [3:0]     OE_DATA_110_const_net_16;
wire   [3:0]     OE_DATA_111_const_net_16;
wire   [3:0]     OE_DATA_112_const_net_16;
wire   [3:0]     OE_DATA_113_const_net_16;
wire   [3:0]     OE_DATA_114_const_net_16;
wire   [3:0]     OE_DATA_115_const_net_16;
wire   [3:0]     OE_DATA_116_const_net_16;
wire   [3:0]     OE_DATA_117_const_net_16;
wire   [3:0]     OE_DATA_118_const_net_16;
wire   [3:0]     OE_DATA_119_const_net_16;
wire   [3:0]     OE_DATA_120_const_net_16;
wire   [3:0]     OE_DATA_121_const_net_16;
wire   [3:0]     OE_DATA_122_const_net_16;
wire   [3:0]     OE_DATA_123_const_net_16;
wire   [3:0]     OE_DATA_124_const_net_16;
wire   [3:0]     OE_DATA_125_const_net_16;
wire   [3:0]     OE_DATA_126_const_net_16;
wire   [3:0]     OE_DATA_127_const_net_16;
wire   [7:0]     PAD_I_const_net_3;
wire   [7:0]     PAD_N_const_net_3;
wire   [7:0]     PAD_I_N_const_net_3;
wire   [7:0]     TX_DATA_1_const_net_13;
wire   [7:0]     TX_DATA_2_const_net_15;
wire   [7:0]     TX_DATA_3_const_net_15;
wire   [7:0]     TX_DATA_4_const_net_15;
wire   [7:0]     TX_DATA_5_const_net_15;
wire   [7:0]     TX_DATA_6_const_net_15;
wire   [7:0]     TX_DATA_7_const_net_15;
wire   [7:0]     TX_DATA_8_const_net_16;
wire   [7:0]     TX_DATA_9_const_net_16;
wire   [7:0]     TX_DATA_10_const_net_16;
wire   [7:0]     TX_DATA_11_const_net_16;
wire   [7:0]     TX_DATA_12_const_net_17;
wire   [7:0]     TX_DATA_13_const_net_17;
wire   [7:0]     TX_DATA_14_const_net_17;
wire   [7:0]     TX_DATA_15_const_net_17;
wire   [7:0]     TX_DATA_16_const_net_17;
wire   [7:0]     TX_DATA_17_const_net_17;
wire   [7:0]     TX_DATA_18_const_net_17;
wire   [7:0]     TX_DATA_19_const_net_17;
wire   [7:0]     TX_DATA_20_const_net_17;
wire   [7:0]     TX_DATA_21_const_net_17;
wire   [7:0]     TX_DATA_22_const_net_17;
wire   [7:0]     TX_DATA_23_const_net_17;
wire   [7:0]     TX_DATA_24_const_net_17;
wire   [7:0]     TX_DATA_25_const_net_17;
wire   [7:0]     TX_DATA_26_const_net_17;
wire   [7:0]     TX_DATA_27_const_net_17;
wire   [7:0]     TX_DATA_28_const_net_17;
wire   [7:0]     TX_DATA_29_const_net_17;
wire   [7:0]     TX_DATA_30_const_net_17;
wire   [7:0]     TX_DATA_31_const_net_17;
wire   [7:0]     TX_DATA_32_const_net_17;
wire   [7:0]     TX_DATA_33_const_net_17;
wire   [7:0]     TX_DATA_34_const_net_17;
wire   [7:0]     TX_DATA_35_const_net_17;
wire   [7:0]     TX_DATA_36_const_net_17;
wire   [7:0]     TX_DATA_37_const_net_17;
wire   [7:0]     TX_DATA_38_const_net_17;
wire   [7:0]     TX_DATA_39_const_net_17;
wire   [7:0]     TX_DATA_40_const_net_17;
wire   [7:0]     TX_DATA_41_const_net_17;
wire   [7:0]     TX_DATA_42_const_net_17;
wire   [7:0]     TX_DATA_43_const_net_17;
wire   [7:0]     TX_DATA_44_const_net_17;
wire   [7:0]     TX_DATA_45_const_net_17;
wire   [7:0]     TX_DATA_46_const_net_17;
wire   [7:0]     TX_DATA_47_const_net_17;
wire   [7:0]     TX_DATA_48_const_net_17;
wire   [7:0]     TX_DATA_49_const_net_17;
wire   [7:0]     TX_DATA_50_const_net_17;
wire   [7:0]     TX_DATA_51_const_net_17;
wire   [7:0]     TX_DATA_52_const_net_17;
wire   [7:0]     TX_DATA_53_const_net_17;
wire   [7:0]     TX_DATA_54_const_net_17;
wire   [7:0]     TX_DATA_55_const_net_17;
wire   [7:0]     TX_DATA_56_const_net_17;
wire   [7:0]     TX_DATA_57_const_net_17;
wire   [7:0]     TX_DATA_58_const_net_17;
wire   [7:0]     TX_DATA_59_const_net_17;
wire   [7:0]     TX_DATA_60_const_net_17;
wire   [7:0]     TX_DATA_61_const_net_17;
wire   [7:0]     TX_DATA_62_const_net_17;
wire   [7:0]     TX_DATA_63_const_net_17;
wire   [7:0]     TX_DATA_64_const_net_17;
wire   [7:0]     TX_DATA_65_const_net_17;
wire   [7:0]     TX_DATA_66_const_net_17;
wire   [7:0]     TX_DATA_67_const_net_17;
wire   [7:0]     TX_DATA_68_const_net_17;
wire   [7:0]     TX_DATA_69_const_net_17;
wire   [7:0]     TX_DATA_70_const_net_17;
wire   [7:0]     TX_DATA_71_const_net_17;
wire   [7:0]     TX_DATA_72_const_net_17;
wire   [7:0]     TX_DATA_73_const_net_17;
wire   [7:0]     TX_DATA_74_const_net_17;
wire   [7:0]     TX_DATA_75_const_net_17;
wire   [7:0]     TX_DATA_76_const_net_17;
wire   [7:0]     TX_DATA_77_const_net_17;
wire   [7:0]     TX_DATA_78_const_net_17;
wire   [7:0]     TX_DATA_79_const_net_17;
wire   [7:0]     TX_DATA_80_const_net_17;
wire   [7:0]     TX_DATA_81_const_net_17;
wire   [7:0]     TX_DATA_82_const_net_17;
wire   [7:0]     TX_DATA_83_const_net_17;
wire   [7:0]     TX_DATA_84_const_net_17;
wire   [7:0]     TX_DATA_85_const_net_17;
wire   [7:0]     TX_DATA_86_const_net_17;
wire   [7:0]     TX_DATA_87_const_net_17;
wire   [7:0]     TX_DATA_88_const_net_17;
wire   [7:0]     TX_DATA_89_const_net_17;
wire   [7:0]     TX_DATA_90_const_net_17;
wire   [7:0]     TX_DATA_91_const_net_17;
wire   [7:0]     TX_DATA_92_const_net_17;
wire   [7:0]     TX_DATA_93_const_net_17;
wire   [7:0]     TX_DATA_94_const_net_17;
wire   [7:0]     TX_DATA_95_const_net_17;
wire   [7:0]     TX_DATA_96_const_net_17;
wire   [7:0]     TX_DATA_97_const_net_17;
wire   [7:0]     TX_DATA_98_const_net_17;
wire   [7:0]     TX_DATA_99_const_net_17;
wire   [7:0]     TX_DATA_100_const_net_17;
wire   [7:0]     TX_DATA_101_const_net_17;
wire   [7:0]     TX_DATA_102_const_net_17;
wire   [7:0]     TX_DATA_103_const_net_17;
wire   [7:0]     TX_DATA_104_const_net_17;
wire   [7:0]     TX_DATA_105_const_net_17;
wire   [7:0]     TX_DATA_106_const_net_17;
wire   [7:0]     TX_DATA_107_const_net_17;
wire   [7:0]     TX_DATA_108_const_net_17;
wire   [7:0]     TX_DATA_109_const_net_17;
wire   [7:0]     TX_DATA_110_const_net_17;
wire   [7:0]     TX_DATA_111_const_net_17;
wire   [7:0]     TX_DATA_112_const_net_17;
wire   [7:0]     TX_DATA_113_const_net_17;
wire   [7:0]     TX_DATA_114_const_net_17;
wire   [7:0]     TX_DATA_115_const_net_17;
wire   [7:0]     TX_DATA_116_const_net_17;
wire   [7:0]     TX_DATA_117_const_net_17;
wire   [7:0]     TX_DATA_118_const_net_17;
wire   [7:0]     TX_DATA_119_const_net_17;
wire   [7:0]     TX_DATA_120_const_net_17;
wire   [7:0]     TX_DATA_121_const_net_17;
wire   [7:0]     TX_DATA_122_const_net_17;
wire   [7:0]     TX_DATA_123_const_net_17;
wire   [7:0]     TX_DATA_124_const_net_17;
wire   [7:0]     TX_DATA_125_const_net_17;
wire   [7:0]     TX_DATA_126_const_net_17;
wire   [7:0]     TX_DATA_127_const_net_17;
wire   [3:0]     OE_DATA_1_const_net_16;
wire   [3:0]     OE_DATA_2_const_net_16;
wire   [3:0]     OE_DATA_3_const_net_16;
wire   [3:0]     OE_DATA_4_const_net_16;
wire   [3:0]     OE_DATA_5_const_net_16;
wire   [3:0]     OE_DATA_6_const_net_16;
wire   [3:0]     OE_DATA_7_const_net_16;
wire   [3:0]     OE_DATA_8_const_net_17;
wire   [3:0]     OE_DATA_9_const_net_17;
wire   [3:0]     OE_DATA_10_const_net_17;
wire   [3:0]     OE_DATA_11_const_net_17;
wire   [3:0]     OE_DATA_12_const_net_17;
wire   [3:0]     OE_DATA_13_const_net_17;
wire   [3:0]     OE_DATA_14_const_net_17;
wire   [3:0]     OE_DATA_15_const_net_17;
wire   [3:0]     OE_DATA_16_const_net_17;
wire   [3:0]     OE_DATA_17_const_net_17;
wire   [3:0]     OE_DATA_18_const_net_17;
wire   [3:0]     OE_DATA_19_const_net_17;
wire   [3:0]     OE_DATA_20_const_net_17;
wire   [3:0]     OE_DATA_21_const_net_17;
wire   [3:0]     OE_DATA_22_const_net_17;
wire   [3:0]     OE_DATA_23_const_net_17;
wire   [3:0]     OE_DATA_24_const_net_17;
wire   [3:0]     OE_DATA_25_const_net_17;
wire   [3:0]     OE_DATA_26_const_net_17;
wire   [3:0]     OE_DATA_27_const_net_17;
wire   [3:0]     OE_DATA_28_const_net_17;
wire   [3:0]     OE_DATA_29_const_net_17;
wire   [3:0]     OE_DATA_30_const_net_17;
wire   [3:0]     OE_DATA_31_const_net_17;
wire   [3:0]     OE_DATA_32_const_net_17;
wire   [3:0]     OE_DATA_33_const_net_17;
wire   [3:0]     OE_DATA_34_const_net_17;
wire   [3:0]     OE_DATA_35_const_net_17;
wire   [3:0]     OE_DATA_36_const_net_17;
wire   [3:0]     OE_DATA_37_const_net_17;
wire   [3:0]     OE_DATA_38_const_net_17;
wire   [3:0]     OE_DATA_39_const_net_17;
wire   [3:0]     OE_DATA_40_const_net_17;
wire   [3:0]     OE_DATA_41_const_net_17;
wire   [3:0]     OE_DATA_42_const_net_17;
wire   [3:0]     OE_DATA_43_const_net_17;
wire   [3:0]     OE_DATA_44_const_net_17;
wire   [3:0]     OE_DATA_45_const_net_17;
wire   [3:0]     OE_DATA_46_const_net_17;
wire   [3:0]     OE_DATA_47_const_net_17;
wire   [3:0]     OE_DATA_48_const_net_17;
wire   [3:0]     OE_DATA_49_const_net_17;
wire   [3:0]     OE_DATA_50_const_net_17;
wire   [3:0]     OE_DATA_51_const_net_17;
wire   [3:0]     OE_DATA_52_const_net_17;
wire   [3:0]     OE_DATA_53_const_net_17;
wire   [3:0]     OE_DATA_54_const_net_17;
wire   [3:0]     OE_DATA_55_const_net_17;
wire   [3:0]     OE_DATA_56_const_net_17;
wire   [3:0]     OE_DATA_57_const_net_17;
wire   [3:0]     OE_DATA_58_const_net_17;
wire   [3:0]     OE_DATA_59_const_net_17;
wire   [3:0]     OE_DATA_60_const_net_17;
wire   [3:0]     OE_DATA_61_const_net_17;
wire   [3:0]     OE_DATA_62_const_net_17;
wire   [3:0]     OE_DATA_63_const_net_17;
wire   [3:0]     OE_DATA_64_const_net_17;
wire   [3:0]     OE_DATA_65_const_net_17;
wire   [3:0]     OE_DATA_66_const_net_17;
wire   [3:0]     OE_DATA_67_const_net_17;
wire   [3:0]     OE_DATA_68_const_net_17;
wire   [3:0]     OE_DATA_69_const_net_17;
wire   [3:0]     OE_DATA_70_const_net_17;
wire   [3:0]     OE_DATA_71_const_net_17;
wire   [3:0]     OE_DATA_72_const_net_17;
wire   [3:0]     OE_DATA_73_const_net_17;
wire   [3:0]     OE_DATA_74_const_net_17;
wire   [3:0]     OE_DATA_75_const_net_17;
wire   [3:0]     OE_DATA_76_const_net_17;
wire   [3:0]     OE_DATA_77_const_net_17;
wire   [3:0]     OE_DATA_78_const_net_17;
wire   [3:0]     OE_DATA_79_const_net_17;
wire   [3:0]     OE_DATA_80_const_net_17;
wire   [3:0]     OE_DATA_81_const_net_17;
wire   [3:0]     OE_DATA_82_const_net_17;
wire   [3:0]     OE_DATA_83_const_net_17;
wire   [3:0]     OE_DATA_84_const_net_17;
wire   [3:0]     OE_DATA_85_const_net_17;
wire   [3:0]     OE_DATA_86_const_net_17;
wire   [3:0]     OE_DATA_87_const_net_17;
wire   [3:0]     OE_DATA_88_const_net_17;
wire   [3:0]     OE_DATA_89_const_net_17;
wire   [3:0]     OE_DATA_90_const_net_17;
wire   [3:0]     OE_DATA_91_const_net_17;
wire   [3:0]     OE_DATA_92_const_net_17;
wire   [3:0]     OE_DATA_93_const_net_17;
wire   [3:0]     OE_DATA_94_const_net_17;
wire   [3:0]     OE_DATA_95_const_net_17;
wire   [3:0]     OE_DATA_96_const_net_17;
wire   [3:0]     OE_DATA_97_const_net_17;
wire   [3:0]     OE_DATA_98_const_net_17;
wire   [3:0]     OE_DATA_99_const_net_17;
wire   [3:0]     OE_DATA_100_const_net_17;
wire   [3:0]     OE_DATA_101_const_net_17;
wire   [3:0]     OE_DATA_102_const_net_17;
wire   [3:0]     OE_DATA_103_const_net_17;
wire   [3:0]     OE_DATA_104_const_net_17;
wire   [3:0]     OE_DATA_105_const_net_17;
wire   [3:0]     OE_DATA_106_const_net_17;
wire   [3:0]     OE_DATA_107_const_net_17;
wire   [3:0]     OE_DATA_108_const_net_17;
wire   [3:0]     OE_DATA_109_const_net_17;
wire   [3:0]     OE_DATA_110_const_net_17;
wire   [3:0]     OE_DATA_111_const_net_17;
wire   [3:0]     OE_DATA_112_const_net_17;
wire   [3:0]     OE_DATA_113_const_net_17;
wire   [3:0]     OE_DATA_114_const_net_17;
wire   [3:0]     OE_DATA_115_const_net_17;
wire   [3:0]     OE_DATA_116_const_net_17;
wire   [3:0]     OE_DATA_117_const_net_17;
wire   [3:0]     OE_DATA_118_const_net_17;
wire   [3:0]     OE_DATA_119_const_net_17;
wire   [3:0]     OE_DATA_120_const_net_17;
wire   [3:0]     OE_DATA_121_const_net_17;
wire   [3:0]     OE_DATA_122_const_net_17;
wire   [3:0]     OE_DATA_123_const_net_17;
wire   [3:0]     OE_DATA_124_const_net_17;
wire   [3:0]     OE_DATA_125_const_net_17;
wire   [3:0]     OE_DATA_126_const_net_17;
wire   [3:0]     OE_DATA_127_const_net_17;
wire   [1:0]     RX_DQS_90_const_net_15;
wire   [2:0]     FIFO_WR_PTR_const_net_16;
wire   [2:0]     FIFO_RD_PTR_const_net_16;
wire   [2:0]     EYE_MONITOR_LANE_WIDTH_const_net_16;
wire   [1:0]     TX_DATA_1_const_net_14;
wire   [1:0]     TX_DATA_2_const_net_16;
wire   [1:0]     TX_DATA_3_const_net_16;
wire   [1:0]     TX_DATA_4_const_net_16;
wire   [1:0]     TX_DATA_5_const_net_16;
wire   [1:0]     TX_DATA_6_const_net_16;
wire   [1:0]     TX_DATA_7_const_net_16;
wire   [1:0]     TX_DATA_8_const_net_17;
wire   [1:0]     TX_DATA_9_const_net_17;
wire   [1:0]     TX_DATA_10_const_net_17;
wire   [1:0]     TX_DATA_11_const_net_17;
wire   [1:0]     TX_DATA_12_const_net_18;
wire   [1:0]     TX_DATA_13_const_net_18;
wire   [1:0]     TX_DATA_14_const_net_18;
wire   [1:0]     TX_DATA_15_const_net_18;
wire   [1:0]     TX_DATA_16_const_net_18;
wire   [1:0]     TX_DATA_17_const_net_18;
wire   [1:0]     TX_DATA_18_const_net_18;
wire   [1:0]     TX_DATA_19_const_net_18;
wire   [1:0]     TX_DATA_20_const_net_18;
wire   [1:0]     TX_DATA_21_const_net_18;
wire   [1:0]     TX_DATA_22_const_net_18;
wire   [1:0]     TX_DATA_23_const_net_18;
wire   [1:0]     TX_DATA_24_const_net_18;
wire   [1:0]     TX_DATA_25_const_net_18;
wire   [1:0]     TX_DATA_26_const_net_18;
wire   [1:0]     TX_DATA_27_const_net_18;
wire   [1:0]     TX_DATA_28_const_net_18;
wire   [1:0]     TX_DATA_29_const_net_18;
wire   [1:0]     TX_DATA_30_const_net_18;
wire   [1:0]     TX_DATA_31_const_net_18;
wire   [1:0]     TX_DATA_32_const_net_18;
wire   [1:0]     TX_DATA_33_const_net_18;
wire   [1:0]     TX_DATA_34_const_net_18;
wire   [1:0]     TX_DATA_35_const_net_18;
wire   [1:0]     TX_DATA_36_const_net_18;
wire   [1:0]     TX_DATA_37_const_net_18;
wire   [1:0]     TX_DATA_38_const_net_18;
wire   [1:0]     TX_DATA_39_const_net_18;
wire   [1:0]     TX_DATA_40_const_net_18;
wire   [1:0]     TX_DATA_41_const_net_18;
wire   [1:0]     TX_DATA_42_const_net_18;
wire   [1:0]     TX_DATA_43_const_net_18;
wire   [1:0]     TX_DATA_44_const_net_18;
wire   [1:0]     TX_DATA_45_const_net_18;
wire   [1:0]     TX_DATA_46_const_net_18;
wire   [1:0]     TX_DATA_47_const_net_18;
wire   [1:0]     TX_DATA_48_const_net_18;
wire   [1:0]     TX_DATA_49_const_net_18;
wire   [1:0]     TX_DATA_50_const_net_18;
wire   [1:0]     TX_DATA_51_const_net_18;
wire   [1:0]     TX_DATA_52_const_net_18;
wire   [1:0]     TX_DATA_53_const_net_18;
wire   [1:0]     TX_DATA_54_const_net_18;
wire   [1:0]     TX_DATA_55_const_net_18;
wire   [1:0]     TX_DATA_56_const_net_18;
wire   [1:0]     TX_DATA_57_const_net_18;
wire   [1:0]     TX_DATA_58_const_net_18;
wire   [1:0]     TX_DATA_59_const_net_18;
wire   [1:0]     TX_DATA_60_const_net_18;
wire   [1:0]     TX_DATA_61_const_net_18;
wire   [1:0]     TX_DATA_62_const_net_18;
wire   [1:0]     TX_DATA_63_const_net_18;
wire   [1:0]     TX_DATA_64_const_net_18;
wire   [1:0]     TX_DATA_65_const_net_18;
wire   [1:0]     TX_DATA_66_const_net_18;
wire   [1:0]     TX_DATA_67_const_net_18;
wire   [1:0]     TX_DATA_68_const_net_18;
wire   [1:0]     TX_DATA_69_const_net_18;
wire   [1:0]     TX_DATA_70_const_net_18;
wire   [1:0]     TX_DATA_71_const_net_18;
wire   [1:0]     TX_DATA_72_const_net_18;
wire   [1:0]     TX_DATA_73_const_net_18;
wire   [1:0]     TX_DATA_74_const_net_18;
wire   [1:0]     TX_DATA_75_const_net_18;
wire   [1:0]     TX_DATA_76_const_net_18;
wire   [1:0]     TX_DATA_77_const_net_18;
wire   [1:0]     TX_DATA_78_const_net_18;
wire   [1:0]     TX_DATA_79_const_net_18;
wire   [1:0]     TX_DATA_80_const_net_18;
wire   [1:0]     TX_DATA_81_const_net_18;
wire   [1:0]     TX_DATA_82_const_net_18;
wire   [1:0]     TX_DATA_83_const_net_18;
wire   [1:0]     TX_DATA_84_const_net_18;
wire   [1:0]     TX_DATA_85_const_net_18;
wire   [1:0]     TX_DATA_86_const_net_18;
wire   [1:0]     TX_DATA_87_const_net_18;
wire   [1:0]     TX_DATA_88_const_net_18;
wire   [1:0]     TX_DATA_89_const_net_18;
wire   [1:0]     TX_DATA_90_const_net_18;
wire   [1:0]     TX_DATA_91_const_net_18;
wire   [1:0]     TX_DATA_92_const_net_18;
wire   [1:0]     TX_DATA_93_const_net_18;
wire   [1:0]     TX_DATA_94_const_net_18;
wire   [1:0]     TX_DATA_95_const_net_18;
wire   [1:0]     TX_DATA_96_const_net_18;
wire   [1:0]     TX_DATA_97_const_net_18;
wire   [1:0]     TX_DATA_98_const_net_18;
wire   [1:0]     TX_DATA_99_const_net_18;
wire   [1:0]     TX_DATA_100_const_net_18;
wire   [1:0]     TX_DATA_101_const_net_18;
wire   [1:0]     TX_DATA_102_const_net_18;
wire   [1:0]     TX_DATA_103_const_net_18;
wire   [1:0]     TX_DATA_104_const_net_18;
wire   [1:0]     TX_DATA_105_const_net_18;
wire   [1:0]     TX_DATA_106_const_net_18;
wire   [1:0]     TX_DATA_107_const_net_18;
wire   [1:0]     TX_DATA_108_const_net_18;
wire   [1:0]     TX_DATA_109_const_net_18;
wire   [1:0]     TX_DATA_110_const_net_18;
wire   [1:0]     TX_DATA_111_const_net_18;
wire   [1:0]     TX_DATA_112_const_net_18;
wire   [1:0]     TX_DATA_113_const_net_18;
wire   [1:0]     TX_DATA_114_const_net_18;
wire   [1:0]     TX_DATA_115_const_net_18;
wire   [1:0]     TX_DATA_116_const_net_18;
wire   [1:0]     TX_DATA_117_const_net_18;
wire   [1:0]     TX_DATA_118_const_net_18;
wire   [1:0]     TX_DATA_119_const_net_18;
wire   [1:0]     TX_DATA_120_const_net_18;
wire   [1:0]     TX_DATA_121_const_net_18;
wire   [1:0]     TX_DATA_122_const_net_18;
wire   [1:0]     TX_DATA_123_const_net_18;
wire   [1:0]     TX_DATA_124_const_net_18;
wire   [1:0]     TX_DATA_125_const_net_18;
wire   [1:0]     TX_DATA_126_const_net_18;
wire   [1:0]     TX_DATA_127_const_net_18;
wire   [1:0]     OE_DATA_1_const_net_17;
wire   [1:0]     OE_DATA_2_const_net_17;
wire   [1:0]     OE_DATA_3_const_net_17;
wire   [1:0]     OE_DATA_4_const_net_17;
wire   [1:0]     OE_DATA_5_const_net_17;
wire   [1:0]     OE_DATA_6_const_net_17;
wire   [1:0]     OE_DATA_7_const_net_17;
wire   [1:0]     OE_DATA_8_const_net_18;
wire   [1:0]     OE_DATA_9_const_net_18;
wire   [1:0]     OE_DATA_10_const_net_18;
wire   [1:0]     OE_DATA_11_const_net_18;
wire   [1:0]     OE_DATA_12_const_net_18;
wire   [1:0]     OE_DATA_13_const_net_18;
wire   [1:0]     OE_DATA_14_const_net_18;
wire   [1:0]     OE_DATA_15_const_net_18;
wire   [1:0]     OE_DATA_16_const_net_18;
wire   [1:0]     OE_DATA_17_const_net_18;
wire   [1:0]     OE_DATA_18_const_net_18;
wire   [1:0]     OE_DATA_19_const_net_18;
wire   [1:0]     OE_DATA_20_const_net_18;
wire   [1:0]     OE_DATA_21_const_net_18;
wire   [1:0]     OE_DATA_22_const_net_18;
wire   [1:0]     OE_DATA_23_const_net_18;
wire   [1:0]     OE_DATA_24_const_net_18;
wire   [1:0]     OE_DATA_25_const_net_18;
wire   [1:0]     OE_DATA_26_const_net_18;
wire   [1:0]     OE_DATA_27_const_net_18;
wire   [1:0]     OE_DATA_28_const_net_18;
wire   [1:0]     OE_DATA_29_const_net_18;
wire   [1:0]     OE_DATA_30_const_net_18;
wire   [1:0]     OE_DATA_31_const_net_18;
wire   [1:0]     OE_DATA_32_const_net_18;
wire   [1:0]     OE_DATA_33_const_net_18;
wire   [1:0]     OE_DATA_34_const_net_18;
wire   [1:0]     OE_DATA_35_const_net_18;
wire   [1:0]     OE_DATA_36_const_net_18;
wire   [1:0]     OE_DATA_37_const_net_18;
wire   [1:0]     OE_DATA_38_const_net_18;
wire   [1:0]     OE_DATA_39_const_net_18;
wire   [1:0]     OE_DATA_40_const_net_18;
wire   [1:0]     OE_DATA_41_const_net_18;
wire   [1:0]     OE_DATA_42_const_net_18;
wire   [1:0]     OE_DATA_43_const_net_18;
wire   [1:0]     OE_DATA_44_const_net_18;
wire   [1:0]     OE_DATA_45_const_net_18;
wire   [1:0]     OE_DATA_46_const_net_18;
wire   [1:0]     OE_DATA_47_const_net_18;
wire   [1:0]     OE_DATA_48_const_net_18;
wire   [1:0]     OE_DATA_49_const_net_18;
wire   [1:0]     OE_DATA_50_const_net_18;
wire   [1:0]     OE_DATA_51_const_net_18;
wire   [1:0]     OE_DATA_52_const_net_18;
wire   [1:0]     OE_DATA_53_const_net_18;
wire   [1:0]     OE_DATA_54_const_net_18;
wire   [1:0]     OE_DATA_55_const_net_18;
wire   [1:0]     OE_DATA_56_const_net_18;
wire   [1:0]     OE_DATA_57_const_net_18;
wire   [1:0]     OE_DATA_58_const_net_18;
wire   [1:0]     OE_DATA_59_const_net_18;
wire   [1:0]     OE_DATA_60_const_net_18;
wire   [1:0]     OE_DATA_61_const_net_18;
wire   [1:0]     OE_DATA_62_const_net_18;
wire   [1:0]     OE_DATA_63_const_net_18;
wire   [1:0]     OE_DATA_64_const_net_18;
wire   [1:0]     OE_DATA_65_const_net_18;
wire   [1:0]     OE_DATA_66_const_net_18;
wire   [1:0]     OE_DATA_67_const_net_18;
wire   [1:0]     OE_DATA_68_const_net_18;
wire   [1:0]     OE_DATA_69_const_net_18;
wire   [1:0]     OE_DATA_70_const_net_18;
wire   [1:0]     OE_DATA_71_const_net_18;
wire   [1:0]     OE_DATA_72_const_net_18;
wire   [1:0]     OE_DATA_73_const_net_18;
wire   [1:0]     OE_DATA_74_const_net_18;
wire   [1:0]     OE_DATA_75_const_net_18;
wire   [1:0]     OE_DATA_76_const_net_18;
wire   [1:0]     OE_DATA_77_const_net_18;
wire   [1:0]     OE_DATA_78_const_net_18;
wire   [1:0]     OE_DATA_79_const_net_18;
wire   [1:0]     OE_DATA_80_const_net_18;
wire   [1:0]     OE_DATA_81_const_net_18;
wire   [1:0]     OE_DATA_82_const_net_18;
wire   [1:0]     OE_DATA_83_const_net_18;
wire   [1:0]     OE_DATA_84_const_net_18;
wire   [1:0]     OE_DATA_85_const_net_18;
wire   [1:0]     OE_DATA_86_const_net_18;
wire   [1:0]     OE_DATA_87_const_net_18;
wire   [1:0]     OE_DATA_88_const_net_18;
wire   [1:0]     OE_DATA_89_const_net_18;
wire   [1:0]     OE_DATA_90_const_net_18;
wire   [1:0]     OE_DATA_91_const_net_18;
wire   [1:0]     OE_DATA_92_const_net_18;
wire   [1:0]     OE_DATA_93_const_net_18;
wire   [1:0]     OE_DATA_94_const_net_18;
wire   [1:0]     OE_DATA_95_const_net_18;
wire   [1:0]     OE_DATA_96_const_net_18;
wire   [1:0]     OE_DATA_97_const_net_18;
wire   [1:0]     OE_DATA_98_const_net_18;
wire   [1:0]     OE_DATA_99_const_net_18;
wire   [1:0]     OE_DATA_100_const_net_18;
wire   [1:0]     OE_DATA_101_const_net_18;
wire   [1:0]     OE_DATA_102_const_net_18;
wire   [1:0]     OE_DATA_103_const_net_18;
wire   [1:0]     OE_DATA_104_const_net_18;
wire   [1:0]     OE_DATA_105_const_net_18;
wire   [1:0]     OE_DATA_106_const_net_18;
wire   [1:0]     OE_DATA_107_const_net_18;
wire   [1:0]     OE_DATA_108_const_net_18;
wire   [1:0]     OE_DATA_109_const_net_18;
wire   [1:0]     OE_DATA_110_const_net_18;
wire   [1:0]     OE_DATA_111_const_net_18;
wire   [1:0]     OE_DATA_112_const_net_18;
wire   [1:0]     OE_DATA_113_const_net_18;
wire   [1:0]     OE_DATA_114_const_net_18;
wire   [1:0]     OE_DATA_115_const_net_18;
wire   [1:0]     OE_DATA_116_const_net_18;
wire   [1:0]     OE_DATA_117_const_net_18;
wire   [1:0]     OE_DATA_118_const_net_18;
wire   [1:0]     OE_DATA_119_const_net_18;
wire   [1:0]     OE_DATA_120_const_net_18;
wire   [1:0]     OE_DATA_121_const_net_18;
wire   [1:0]     OE_DATA_122_const_net_18;
wire   [1:0]     OE_DATA_123_const_net_18;
wire   [1:0]     OE_DATA_124_const_net_18;
wire   [1:0]     OE_DATA_125_const_net_18;
wire   [1:0]     OE_DATA_126_const_net_18;
wire   [1:0]     OE_DATA_127_const_net_18;
wire   [1:0]     RX_DQS_90_const_net_16;
wire   [2:0]     EYE_MONITOR_LANE_WIDTH_const_net_17;
wire   [7:0]     TX_DATA_1_const_net_15;
wire   [7:0]     TX_DATA_2_const_net_17;
wire   [7:0]     TX_DATA_3_const_net_17;
wire   [7:0]     TX_DATA_4_const_net_17;
wire   [7:0]     TX_DATA_5_const_net_17;
wire   [7:0]     TX_DATA_6_const_net_17;
wire   [7:0]     TX_DATA_7_const_net_17;
wire   [7:0]     TX_DATA_8_const_net_18;
wire   [7:0]     TX_DATA_9_const_net_18;
wire   [7:0]     TX_DATA_10_const_net_18;
wire   [7:0]     TX_DATA_11_const_net_18;
wire   [7:0]     TX_DATA_12_const_net_19;
wire   [7:0]     TX_DATA_13_const_net_19;
wire   [7:0]     TX_DATA_14_const_net_19;
wire   [7:0]     TX_DATA_15_const_net_19;
wire   [7:0]     TX_DATA_16_const_net_19;
wire   [7:0]     TX_DATA_17_const_net_19;
wire   [7:0]     TX_DATA_18_const_net_19;
wire   [7:0]     TX_DATA_19_const_net_19;
wire   [7:0]     TX_DATA_20_const_net_19;
wire   [7:0]     TX_DATA_21_const_net_19;
wire   [7:0]     TX_DATA_22_const_net_19;
wire   [7:0]     TX_DATA_23_const_net_19;
wire   [7:0]     TX_DATA_24_const_net_19;
wire   [7:0]     TX_DATA_25_const_net_19;
wire   [7:0]     TX_DATA_26_const_net_19;
wire   [7:0]     TX_DATA_27_const_net_19;
wire   [7:0]     TX_DATA_28_const_net_19;
wire   [7:0]     TX_DATA_29_const_net_19;
wire   [7:0]     TX_DATA_30_const_net_19;
wire   [7:0]     TX_DATA_31_const_net_19;
wire   [7:0]     TX_DATA_32_const_net_19;
wire   [7:0]     TX_DATA_33_const_net_19;
wire   [7:0]     TX_DATA_34_const_net_19;
wire   [7:0]     TX_DATA_35_const_net_19;
wire   [7:0]     TX_DATA_36_const_net_19;
wire   [7:0]     TX_DATA_37_const_net_19;
wire   [7:0]     TX_DATA_38_const_net_19;
wire   [7:0]     TX_DATA_39_const_net_19;
wire   [7:0]     TX_DATA_40_const_net_19;
wire   [7:0]     TX_DATA_41_const_net_19;
wire   [7:0]     TX_DATA_42_const_net_19;
wire   [7:0]     TX_DATA_43_const_net_19;
wire   [7:0]     TX_DATA_44_const_net_19;
wire   [7:0]     TX_DATA_45_const_net_19;
wire   [7:0]     TX_DATA_46_const_net_19;
wire   [7:0]     TX_DATA_47_const_net_19;
wire   [7:0]     TX_DATA_48_const_net_19;
wire   [7:0]     TX_DATA_49_const_net_19;
wire   [7:0]     TX_DATA_50_const_net_19;
wire   [7:0]     TX_DATA_51_const_net_19;
wire   [7:0]     TX_DATA_52_const_net_19;
wire   [7:0]     TX_DATA_53_const_net_19;
wire   [7:0]     TX_DATA_54_const_net_19;
wire   [7:0]     TX_DATA_55_const_net_19;
wire   [7:0]     TX_DATA_56_const_net_19;
wire   [7:0]     TX_DATA_57_const_net_19;
wire   [7:0]     TX_DATA_58_const_net_19;
wire   [7:0]     TX_DATA_59_const_net_19;
wire   [7:0]     TX_DATA_60_const_net_19;
wire   [7:0]     TX_DATA_61_const_net_19;
wire   [7:0]     TX_DATA_62_const_net_19;
wire   [7:0]     TX_DATA_63_const_net_19;
wire   [7:0]     TX_DATA_64_const_net_19;
wire   [7:0]     TX_DATA_65_const_net_19;
wire   [7:0]     TX_DATA_66_const_net_19;
wire   [7:0]     TX_DATA_67_const_net_19;
wire   [7:0]     TX_DATA_68_const_net_19;
wire   [7:0]     TX_DATA_69_const_net_19;
wire   [7:0]     TX_DATA_70_const_net_19;
wire   [7:0]     TX_DATA_71_const_net_19;
wire   [7:0]     TX_DATA_72_const_net_19;
wire   [7:0]     TX_DATA_73_const_net_19;
wire   [7:0]     TX_DATA_74_const_net_19;
wire   [7:0]     TX_DATA_75_const_net_19;
wire   [7:0]     TX_DATA_76_const_net_19;
wire   [7:0]     TX_DATA_77_const_net_19;
wire   [7:0]     TX_DATA_78_const_net_19;
wire   [7:0]     TX_DATA_79_const_net_19;
wire   [7:0]     TX_DATA_80_const_net_19;
wire   [7:0]     TX_DATA_81_const_net_19;
wire   [7:0]     TX_DATA_82_const_net_19;
wire   [7:0]     TX_DATA_83_const_net_19;
wire   [7:0]     TX_DATA_84_const_net_19;
wire   [7:0]     TX_DATA_85_const_net_19;
wire   [7:0]     TX_DATA_86_const_net_19;
wire   [7:0]     TX_DATA_87_const_net_19;
wire   [7:0]     TX_DATA_88_const_net_19;
wire   [7:0]     TX_DATA_89_const_net_19;
wire   [7:0]     TX_DATA_90_const_net_19;
wire   [7:0]     TX_DATA_91_const_net_19;
wire   [7:0]     TX_DATA_92_const_net_19;
wire   [7:0]     TX_DATA_93_const_net_19;
wire   [7:0]     TX_DATA_94_const_net_19;
wire   [7:0]     TX_DATA_95_const_net_19;
wire   [7:0]     TX_DATA_96_const_net_19;
wire   [7:0]     TX_DATA_97_const_net_19;
wire   [7:0]     TX_DATA_98_const_net_19;
wire   [7:0]     TX_DATA_99_const_net_19;
wire   [7:0]     TX_DATA_100_const_net_19;
wire   [7:0]     TX_DATA_101_const_net_19;
wire   [7:0]     TX_DATA_102_const_net_19;
wire   [7:0]     TX_DATA_103_const_net_19;
wire   [7:0]     TX_DATA_104_const_net_19;
wire   [7:0]     TX_DATA_105_const_net_19;
wire   [7:0]     TX_DATA_106_const_net_19;
wire   [7:0]     TX_DATA_107_const_net_19;
wire   [7:0]     TX_DATA_108_const_net_19;
wire   [7:0]     TX_DATA_109_const_net_19;
wire   [7:0]     TX_DATA_110_const_net_19;
wire   [7:0]     TX_DATA_111_const_net_19;
wire   [7:0]     TX_DATA_112_const_net_19;
wire   [7:0]     TX_DATA_113_const_net_19;
wire   [7:0]     TX_DATA_114_const_net_19;
wire   [7:0]     TX_DATA_115_const_net_19;
wire   [7:0]     TX_DATA_116_const_net_19;
wire   [7:0]     TX_DATA_117_const_net_19;
wire   [7:0]     TX_DATA_118_const_net_19;
wire   [7:0]     TX_DATA_119_const_net_19;
wire   [7:0]     TX_DATA_120_const_net_19;
wire   [7:0]     TX_DATA_121_const_net_19;
wire   [7:0]     TX_DATA_122_const_net_19;
wire   [7:0]     TX_DATA_123_const_net_19;
wire   [7:0]     TX_DATA_124_const_net_19;
wire   [7:0]     TX_DATA_125_const_net_19;
wire   [7:0]     TX_DATA_126_const_net_19;
wire   [7:0]     TX_DATA_127_const_net_19;
wire   [3:0]     OE_DATA_1_const_net_18;
wire   [3:0]     OE_DATA_2_const_net_18;
wire   [3:0]     OE_DATA_3_const_net_18;
wire   [3:0]     OE_DATA_4_const_net_18;
wire   [3:0]     OE_DATA_5_const_net_18;
wire   [3:0]     OE_DATA_6_const_net_18;
wire   [3:0]     OE_DATA_7_const_net_18;
wire   [3:0]     OE_DATA_8_const_net_19;
wire   [3:0]     OE_DATA_9_const_net_19;
wire   [3:0]     OE_DATA_10_const_net_19;
wire   [3:0]     OE_DATA_11_const_net_19;
wire   [3:0]     OE_DATA_12_const_net_19;
wire   [3:0]     OE_DATA_13_const_net_19;
wire   [3:0]     OE_DATA_14_const_net_19;
wire   [3:0]     OE_DATA_15_const_net_19;
wire   [3:0]     OE_DATA_16_const_net_19;
wire   [3:0]     OE_DATA_17_const_net_19;
wire   [3:0]     OE_DATA_18_const_net_19;
wire   [3:0]     OE_DATA_19_const_net_19;
wire   [3:0]     OE_DATA_20_const_net_19;
wire   [3:0]     OE_DATA_21_const_net_19;
wire   [3:0]     OE_DATA_22_const_net_19;
wire   [3:0]     OE_DATA_23_const_net_19;
wire   [3:0]     OE_DATA_24_const_net_19;
wire   [3:0]     OE_DATA_25_const_net_19;
wire   [3:0]     OE_DATA_26_const_net_19;
wire   [3:0]     OE_DATA_27_const_net_19;
wire   [3:0]     OE_DATA_28_const_net_19;
wire   [3:0]     OE_DATA_29_const_net_19;
wire   [3:0]     OE_DATA_30_const_net_19;
wire   [3:0]     OE_DATA_31_const_net_19;
wire   [3:0]     OE_DATA_32_const_net_19;
wire   [3:0]     OE_DATA_33_const_net_19;
wire   [3:0]     OE_DATA_34_const_net_19;
wire   [3:0]     OE_DATA_35_const_net_19;
wire   [3:0]     OE_DATA_36_const_net_19;
wire   [3:0]     OE_DATA_37_const_net_19;
wire   [3:0]     OE_DATA_38_const_net_19;
wire   [3:0]     OE_DATA_39_const_net_19;
wire   [3:0]     OE_DATA_40_const_net_19;
wire   [3:0]     OE_DATA_41_const_net_19;
wire   [3:0]     OE_DATA_42_const_net_19;
wire   [3:0]     OE_DATA_43_const_net_19;
wire   [3:0]     OE_DATA_44_const_net_19;
wire   [3:0]     OE_DATA_45_const_net_19;
wire   [3:0]     OE_DATA_46_const_net_19;
wire   [3:0]     OE_DATA_47_const_net_19;
wire   [3:0]     OE_DATA_48_const_net_19;
wire   [3:0]     OE_DATA_49_const_net_19;
wire   [3:0]     OE_DATA_50_const_net_19;
wire   [3:0]     OE_DATA_51_const_net_19;
wire   [3:0]     OE_DATA_52_const_net_19;
wire   [3:0]     OE_DATA_53_const_net_19;
wire   [3:0]     OE_DATA_54_const_net_19;
wire   [3:0]     OE_DATA_55_const_net_19;
wire   [3:0]     OE_DATA_56_const_net_19;
wire   [3:0]     OE_DATA_57_const_net_19;
wire   [3:0]     OE_DATA_58_const_net_19;
wire   [3:0]     OE_DATA_59_const_net_19;
wire   [3:0]     OE_DATA_60_const_net_19;
wire   [3:0]     OE_DATA_61_const_net_19;
wire   [3:0]     OE_DATA_62_const_net_19;
wire   [3:0]     OE_DATA_63_const_net_19;
wire   [3:0]     OE_DATA_64_const_net_19;
wire   [3:0]     OE_DATA_65_const_net_19;
wire   [3:0]     OE_DATA_66_const_net_19;
wire   [3:0]     OE_DATA_67_const_net_19;
wire   [3:0]     OE_DATA_68_const_net_19;
wire   [3:0]     OE_DATA_69_const_net_19;
wire   [3:0]     OE_DATA_70_const_net_19;
wire   [3:0]     OE_DATA_71_const_net_19;
wire   [3:0]     OE_DATA_72_const_net_19;
wire   [3:0]     OE_DATA_73_const_net_19;
wire   [3:0]     OE_DATA_74_const_net_19;
wire   [3:0]     OE_DATA_75_const_net_19;
wire   [3:0]     OE_DATA_76_const_net_19;
wire   [3:0]     OE_DATA_77_const_net_19;
wire   [3:0]     OE_DATA_78_const_net_19;
wire   [3:0]     OE_DATA_79_const_net_19;
wire   [3:0]     OE_DATA_80_const_net_19;
wire   [3:0]     OE_DATA_81_const_net_19;
wire   [3:0]     OE_DATA_82_const_net_19;
wire   [3:0]     OE_DATA_83_const_net_19;
wire   [3:0]     OE_DATA_84_const_net_19;
wire   [3:0]     OE_DATA_85_const_net_19;
wire   [3:0]     OE_DATA_86_const_net_19;
wire   [3:0]     OE_DATA_87_const_net_19;
wire   [3:0]     OE_DATA_88_const_net_19;
wire   [3:0]     OE_DATA_89_const_net_19;
wire   [3:0]     OE_DATA_90_const_net_19;
wire   [3:0]     OE_DATA_91_const_net_19;
wire   [3:0]     OE_DATA_92_const_net_19;
wire   [3:0]     OE_DATA_93_const_net_19;
wire   [3:0]     OE_DATA_94_const_net_19;
wire   [3:0]     OE_DATA_95_const_net_19;
wire   [3:0]     OE_DATA_96_const_net_19;
wire   [3:0]     OE_DATA_97_const_net_19;
wire   [3:0]     OE_DATA_98_const_net_19;
wire   [3:0]     OE_DATA_99_const_net_19;
wire   [3:0]     OE_DATA_100_const_net_19;
wire   [3:0]     OE_DATA_101_const_net_19;
wire   [3:0]     OE_DATA_102_const_net_19;
wire   [3:0]     OE_DATA_103_const_net_19;
wire   [3:0]     OE_DATA_104_const_net_19;
wire   [3:0]     OE_DATA_105_const_net_19;
wire   [3:0]     OE_DATA_106_const_net_19;
wire   [3:0]     OE_DATA_107_const_net_19;
wire   [3:0]     OE_DATA_108_const_net_19;
wire   [3:0]     OE_DATA_109_const_net_19;
wire   [3:0]     OE_DATA_110_const_net_19;
wire   [3:0]     OE_DATA_111_const_net_19;
wire   [3:0]     OE_DATA_112_const_net_19;
wire   [3:0]     OE_DATA_113_const_net_19;
wire   [3:0]     OE_DATA_114_const_net_19;
wire   [3:0]     OE_DATA_115_const_net_19;
wire   [3:0]     OE_DATA_116_const_net_19;
wire   [3:0]     OE_DATA_117_const_net_19;
wire   [3:0]     OE_DATA_118_const_net_19;
wire   [3:0]     OE_DATA_119_const_net_19;
wire   [3:0]     OE_DATA_120_const_net_19;
wire   [3:0]     OE_DATA_121_const_net_19;
wire   [3:0]     OE_DATA_122_const_net_19;
wire   [3:0]     OE_DATA_123_const_net_19;
wire   [3:0]     OE_DATA_124_const_net_19;
wire   [3:0]     OE_DATA_125_const_net_19;
wire   [3:0]     OE_DATA_126_const_net_19;
wire   [3:0]     OE_DATA_127_const_net_19;
wire   [10:0]    CDR_CLK_B_SEL_const_net_1;
wire   [2:0]     FIFO_WR_PTR_const_net_17;
wire   [2:0]     FIFO_RD_PTR_const_net_17;
wire   [2:0]     EYE_MONITOR_LANE_WIDTH_const_net_18;
wire   [7:0]     TX_DATA_1_const_net_16;
wire   [7:0]     TX_DATA_2_const_net_18;
wire   [7:0]     TX_DATA_3_const_net_18;
wire   [7:0]     TX_DATA_4_const_net_18;
wire   [7:0]     TX_DATA_5_const_net_18;
wire   [7:0]     TX_DATA_6_const_net_18;
wire   [7:0]     TX_DATA_7_const_net_18;
wire   [7:0]     TX_DATA_8_const_net_19;
wire   [7:0]     TX_DATA_9_const_net_19;
wire   [7:0]     TX_DATA_10_const_net_19;
wire   [7:0]     TX_DATA_11_const_net_19;
wire   [7:0]     TX_DATA_12_const_net_20;
wire   [7:0]     TX_DATA_13_const_net_20;
wire   [7:0]     TX_DATA_14_const_net_20;
wire   [7:0]     TX_DATA_15_const_net_20;
wire   [7:0]     TX_DATA_16_const_net_20;
wire   [7:0]     TX_DATA_17_const_net_20;
wire   [7:0]     TX_DATA_18_const_net_20;
wire   [7:0]     TX_DATA_19_const_net_20;
wire   [7:0]     TX_DATA_20_const_net_20;
wire   [7:0]     TX_DATA_21_const_net_20;
wire   [7:0]     TX_DATA_22_const_net_20;
wire   [7:0]     TX_DATA_23_const_net_20;
wire   [7:0]     TX_DATA_24_const_net_20;
wire   [7:0]     TX_DATA_25_const_net_20;
wire   [7:0]     TX_DATA_26_const_net_20;
wire   [7:0]     TX_DATA_27_const_net_20;
wire   [7:0]     TX_DATA_28_const_net_20;
wire   [7:0]     TX_DATA_29_const_net_20;
wire   [7:0]     TX_DATA_30_const_net_20;
wire   [7:0]     TX_DATA_31_const_net_20;
wire   [7:0]     TX_DATA_32_const_net_20;
wire   [7:0]     TX_DATA_33_const_net_20;
wire   [7:0]     TX_DATA_34_const_net_20;
wire   [7:0]     TX_DATA_35_const_net_20;
wire   [7:0]     TX_DATA_36_const_net_20;
wire   [7:0]     TX_DATA_37_const_net_20;
wire   [7:0]     TX_DATA_38_const_net_20;
wire   [7:0]     TX_DATA_39_const_net_20;
wire   [7:0]     TX_DATA_40_const_net_20;
wire   [7:0]     TX_DATA_41_const_net_20;
wire   [7:0]     TX_DATA_42_const_net_20;
wire   [7:0]     TX_DATA_43_const_net_20;
wire   [7:0]     TX_DATA_44_const_net_20;
wire   [7:0]     TX_DATA_45_const_net_20;
wire   [7:0]     TX_DATA_46_const_net_20;
wire   [7:0]     TX_DATA_47_const_net_20;
wire   [7:0]     TX_DATA_48_const_net_20;
wire   [7:0]     TX_DATA_49_const_net_20;
wire   [7:0]     TX_DATA_50_const_net_20;
wire   [7:0]     TX_DATA_51_const_net_20;
wire   [7:0]     TX_DATA_52_const_net_20;
wire   [7:0]     TX_DATA_53_const_net_20;
wire   [7:0]     TX_DATA_54_const_net_20;
wire   [7:0]     TX_DATA_55_const_net_20;
wire   [7:0]     TX_DATA_56_const_net_20;
wire   [7:0]     TX_DATA_57_const_net_20;
wire   [7:0]     TX_DATA_58_const_net_20;
wire   [7:0]     TX_DATA_59_const_net_20;
wire   [7:0]     TX_DATA_60_const_net_20;
wire   [7:0]     TX_DATA_61_const_net_20;
wire   [7:0]     TX_DATA_62_const_net_20;
wire   [7:0]     TX_DATA_63_const_net_20;
wire   [7:0]     TX_DATA_64_const_net_20;
wire   [7:0]     TX_DATA_65_const_net_20;
wire   [7:0]     TX_DATA_66_const_net_20;
wire   [7:0]     TX_DATA_67_const_net_20;
wire   [7:0]     TX_DATA_68_const_net_20;
wire   [7:0]     TX_DATA_69_const_net_20;
wire   [7:0]     TX_DATA_70_const_net_20;
wire   [7:0]     TX_DATA_71_const_net_20;
wire   [7:0]     TX_DATA_72_const_net_20;
wire   [7:0]     TX_DATA_73_const_net_20;
wire   [7:0]     TX_DATA_74_const_net_20;
wire   [7:0]     TX_DATA_75_const_net_20;
wire   [7:0]     TX_DATA_76_const_net_20;
wire   [7:0]     TX_DATA_77_const_net_20;
wire   [7:0]     TX_DATA_78_const_net_20;
wire   [7:0]     TX_DATA_79_const_net_20;
wire   [7:0]     TX_DATA_80_const_net_20;
wire   [7:0]     TX_DATA_81_const_net_20;
wire   [7:0]     TX_DATA_82_const_net_20;
wire   [7:0]     TX_DATA_83_const_net_20;
wire   [7:0]     TX_DATA_84_const_net_20;
wire   [7:0]     TX_DATA_85_const_net_20;
wire   [7:0]     TX_DATA_86_const_net_20;
wire   [7:0]     TX_DATA_87_const_net_20;
wire   [7:0]     TX_DATA_88_const_net_20;
wire   [7:0]     TX_DATA_89_const_net_20;
wire   [7:0]     TX_DATA_90_const_net_20;
wire   [7:0]     TX_DATA_91_const_net_20;
wire   [7:0]     TX_DATA_92_const_net_20;
wire   [7:0]     TX_DATA_93_const_net_20;
wire   [7:0]     TX_DATA_94_const_net_20;
wire   [7:0]     TX_DATA_95_const_net_20;
wire   [7:0]     TX_DATA_96_const_net_20;
wire   [7:0]     TX_DATA_97_const_net_20;
wire   [7:0]     TX_DATA_98_const_net_20;
wire   [7:0]     TX_DATA_99_const_net_20;
wire   [7:0]     TX_DATA_100_const_net_20;
wire   [7:0]     TX_DATA_101_const_net_20;
wire   [7:0]     TX_DATA_102_const_net_20;
wire   [7:0]     TX_DATA_103_const_net_20;
wire   [7:0]     TX_DATA_104_const_net_20;
wire   [7:0]     TX_DATA_105_const_net_20;
wire   [7:0]     TX_DATA_106_const_net_20;
wire   [7:0]     TX_DATA_107_const_net_20;
wire   [7:0]     TX_DATA_108_const_net_20;
wire   [7:0]     TX_DATA_109_const_net_20;
wire   [7:0]     TX_DATA_110_const_net_20;
wire   [7:0]     TX_DATA_111_const_net_20;
wire   [7:0]     TX_DATA_112_const_net_20;
wire   [7:0]     TX_DATA_113_const_net_20;
wire   [7:0]     TX_DATA_114_const_net_20;
wire   [7:0]     TX_DATA_115_const_net_20;
wire   [7:0]     TX_DATA_116_const_net_20;
wire   [7:0]     TX_DATA_117_const_net_20;
wire   [7:0]     TX_DATA_118_const_net_20;
wire   [7:0]     TX_DATA_119_const_net_20;
wire   [7:0]     TX_DATA_120_const_net_20;
wire   [7:0]     TX_DATA_121_const_net_20;
wire   [7:0]     TX_DATA_122_const_net_20;
wire   [7:0]     TX_DATA_123_const_net_20;
wire   [7:0]     TX_DATA_124_const_net_20;
wire   [7:0]     TX_DATA_125_const_net_20;
wire   [7:0]     TX_DATA_126_const_net_20;
wire   [7:0]     TX_DATA_127_const_net_20;
wire   [3:0]     OE_DATA_1_const_net_19;
wire   [3:0]     OE_DATA_2_const_net_19;
wire   [3:0]     OE_DATA_3_const_net_19;
wire   [3:0]     OE_DATA_4_const_net_19;
wire   [3:0]     OE_DATA_5_const_net_19;
wire   [3:0]     OE_DATA_6_const_net_19;
wire   [3:0]     OE_DATA_7_const_net_19;
wire   [3:0]     OE_DATA_8_const_net_20;
wire   [3:0]     OE_DATA_9_const_net_20;
wire   [3:0]     OE_DATA_10_const_net_20;
wire   [3:0]     OE_DATA_11_const_net_20;
wire   [3:0]     OE_DATA_12_const_net_20;
wire   [3:0]     OE_DATA_13_const_net_20;
wire   [3:0]     OE_DATA_14_const_net_20;
wire   [3:0]     OE_DATA_15_const_net_20;
wire   [3:0]     OE_DATA_16_const_net_20;
wire   [3:0]     OE_DATA_17_const_net_20;
wire   [3:0]     OE_DATA_18_const_net_20;
wire   [3:0]     OE_DATA_19_const_net_20;
wire   [3:0]     OE_DATA_20_const_net_20;
wire   [3:0]     OE_DATA_21_const_net_20;
wire   [3:0]     OE_DATA_22_const_net_20;
wire   [3:0]     OE_DATA_23_const_net_20;
wire   [3:0]     OE_DATA_24_const_net_20;
wire   [3:0]     OE_DATA_25_const_net_20;
wire   [3:0]     OE_DATA_26_const_net_20;
wire   [3:0]     OE_DATA_27_const_net_20;
wire   [3:0]     OE_DATA_28_const_net_20;
wire   [3:0]     OE_DATA_29_const_net_20;
wire   [3:0]     OE_DATA_30_const_net_20;
wire   [3:0]     OE_DATA_31_const_net_20;
wire   [3:0]     OE_DATA_32_const_net_20;
wire   [3:0]     OE_DATA_33_const_net_20;
wire   [3:0]     OE_DATA_34_const_net_20;
wire   [3:0]     OE_DATA_35_const_net_20;
wire   [3:0]     OE_DATA_36_const_net_20;
wire   [3:0]     OE_DATA_37_const_net_20;
wire   [3:0]     OE_DATA_38_const_net_20;
wire   [3:0]     OE_DATA_39_const_net_20;
wire   [3:0]     OE_DATA_40_const_net_20;
wire   [3:0]     OE_DATA_41_const_net_20;
wire   [3:0]     OE_DATA_42_const_net_20;
wire   [3:0]     OE_DATA_43_const_net_20;
wire   [3:0]     OE_DATA_44_const_net_20;
wire   [3:0]     OE_DATA_45_const_net_20;
wire   [3:0]     OE_DATA_46_const_net_20;
wire   [3:0]     OE_DATA_47_const_net_20;
wire   [3:0]     OE_DATA_48_const_net_20;
wire   [3:0]     OE_DATA_49_const_net_20;
wire   [3:0]     OE_DATA_50_const_net_20;
wire   [3:0]     OE_DATA_51_const_net_20;
wire   [3:0]     OE_DATA_52_const_net_20;
wire   [3:0]     OE_DATA_53_const_net_20;
wire   [3:0]     OE_DATA_54_const_net_20;
wire   [3:0]     OE_DATA_55_const_net_20;
wire   [3:0]     OE_DATA_56_const_net_20;
wire   [3:0]     OE_DATA_57_const_net_20;
wire   [3:0]     OE_DATA_58_const_net_20;
wire   [3:0]     OE_DATA_59_const_net_20;
wire   [3:0]     OE_DATA_60_const_net_20;
wire   [3:0]     OE_DATA_61_const_net_20;
wire   [3:0]     OE_DATA_62_const_net_20;
wire   [3:0]     OE_DATA_63_const_net_20;
wire   [3:0]     OE_DATA_64_const_net_20;
wire   [3:0]     OE_DATA_65_const_net_20;
wire   [3:0]     OE_DATA_66_const_net_20;
wire   [3:0]     OE_DATA_67_const_net_20;
wire   [3:0]     OE_DATA_68_const_net_20;
wire   [3:0]     OE_DATA_69_const_net_20;
wire   [3:0]     OE_DATA_70_const_net_20;
wire   [3:0]     OE_DATA_71_const_net_20;
wire   [3:0]     OE_DATA_72_const_net_20;
wire   [3:0]     OE_DATA_73_const_net_20;
wire   [3:0]     OE_DATA_74_const_net_20;
wire   [3:0]     OE_DATA_75_const_net_20;
wire   [3:0]     OE_DATA_76_const_net_20;
wire   [3:0]     OE_DATA_77_const_net_20;
wire   [3:0]     OE_DATA_78_const_net_20;
wire   [3:0]     OE_DATA_79_const_net_20;
wire   [3:0]     OE_DATA_80_const_net_20;
wire   [3:0]     OE_DATA_81_const_net_20;
wire   [3:0]     OE_DATA_82_const_net_20;
wire   [3:0]     OE_DATA_83_const_net_20;
wire   [3:0]     OE_DATA_84_const_net_20;
wire   [3:0]     OE_DATA_85_const_net_20;
wire   [3:0]     OE_DATA_86_const_net_20;
wire   [3:0]     OE_DATA_87_const_net_20;
wire   [3:0]     OE_DATA_88_const_net_20;
wire   [3:0]     OE_DATA_89_const_net_20;
wire   [3:0]     OE_DATA_90_const_net_20;
wire   [3:0]     OE_DATA_91_const_net_20;
wire   [3:0]     OE_DATA_92_const_net_20;
wire   [3:0]     OE_DATA_93_const_net_20;
wire   [3:0]     OE_DATA_94_const_net_20;
wire   [3:0]     OE_DATA_95_const_net_20;
wire   [3:0]     OE_DATA_96_const_net_20;
wire   [3:0]     OE_DATA_97_const_net_20;
wire   [3:0]     OE_DATA_98_const_net_20;
wire   [3:0]     OE_DATA_99_const_net_20;
wire   [3:0]     OE_DATA_100_const_net_20;
wire   [3:0]     OE_DATA_101_const_net_20;
wire   [3:0]     OE_DATA_102_const_net_20;
wire   [3:0]     OE_DATA_103_const_net_20;
wire   [3:0]     OE_DATA_104_const_net_20;
wire   [3:0]     OE_DATA_105_const_net_20;
wire   [3:0]     OE_DATA_106_const_net_20;
wire   [3:0]     OE_DATA_107_const_net_20;
wire   [3:0]     OE_DATA_108_const_net_20;
wire   [3:0]     OE_DATA_109_const_net_20;
wire   [3:0]     OE_DATA_110_const_net_20;
wire   [3:0]     OE_DATA_111_const_net_20;
wire   [3:0]     OE_DATA_112_const_net_20;
wire   [3:0]     OE_DATA_113_const_net_20;
wire   [3:0]     OE_DATA_114_const_net_20;
wire   [3:0]     OE_DATA_115_const_net_20;
wire   [3:0]     OE_DATA_116_const_net_20;
wire   [3:0]     OE_DATA_117_const_net_20;
wire   [3:0]     OE_DATA_118_const_net_20;
wire   [3:0]     OE_DATA_119_const_net_20;
wire   [3:0]     OE_DATA_120_const_net_20;
wire   [3:0]     OE_DATA_121_const_net_20;
wire   [3:0]     OE_DATA_122_const_net_20;
wire   [3:0]     OE_DATA_123_const_net_20;
wire   [3:0]     OE_DATA_124_const_net_20;
wire   [3:0]     OE_DATA_125_const_net_20;
wire   [3:0]     OE_DATA_126_const_net_20;
wire   [3:0]     OE_DATA_127_const_net_20;
wire   [7:0]     TX_DATA_8_const_net_20;
wire   [7:0]     TX_DATA_9_const_net_20;
wire   [7:0]     TX_DATA_10_const_net_20;
wire   [7:0]     TX_DATA_11_const_net_20;
wire   [7:0]     TX_DATA_12_const_net_21;
wire   [7:0]     TX_DATA_13_const_net_21;
wire   [7:0]     TX_DATA_14_const_net_21;
wire   [7:0]     TX_DATA_15_const_net_21;
wire   [7:0]     TX_DATA_16_const_net_21;
wire   [7:0]     TX_DATA_17_const_net_21;
wire   [7:0]     TX_DATA_18_const_net_21;
wire   [7:0]     TX_DATA_19_const_net_21;
wire   [7:0]     TX_DATA_20_const_net_21;
wire   [7:0]     TX_DATA_21_const_net_21;
wire   [7:0]     TX_DATA_22_const_net_21;
wire   [7:0]     TX_DATA_23_const_net_21;
wire   [7:0]     TX_DATA_24_const_net_21;
wire   [7:0]     TX_DATA_25_const_net_21;
wire   [7:0]     TX_DATA_26_const_net_21;
wire   [7:0]     TX_DATA_27_const_net_21;
wire   [7:0]     TX_DATA_28_const_net_21;
wire   [7:0]     TX_DATA_29_const_net_21;
wire   [7:0]     TX_DATA_30_const_net_21;
wire   [7:0]     TX_DATA_31_const_net_21;
wire   [7:0]     TX_DATA_32_const_net_21;
wire   [7:0]     TX_DATA_33_const_net_21;
wire   [7:0]     TX_DATA_34_const_net_21;
wire   [7:0]     TX_DATA_35_const_net_21;
wire   [7:0]     TX_DATA_36_const_net_21;
wire   [7:0]     TX_DATA_37_const_net_21;
wire   [7:0]     TX_DATA_38_const_net_21;
wire   [7:0]     TX_DATA_39_const_net_21;
wire   [7:0]     TX_DATA_40_const_net_21;
wire   [7:0]     TX_DATA_41_const_net_21;
wire   [7:0]     TX_DATA_42_const_net_21;
wire   [7:0]     TX_DATA_43_const_net_21;
wire   [7:0]     TX_DATA_44_const_net_21;
wire   [7:0]     TX_DATA_45_const_net_21;
wire   [7:0]     TX_DATA_46_const_net_21;
wire   [7:0]     TX_DATA_47_const_net_21;
wire   [7:0]     TX_DATA_48_const_net_21;
wire   [7:0]     TX_DATA_49_const_net_21;
wire   [7:0]     TX_DATA_50_const_net_21;
wire   [7:0]     TX_DATA_51_const_net_21;
wire   [7:0]     TX_DATA_52_const_net_21;
wire   [7:0]     TX_DATA_53_const_net_21;
wire   [7:0]     TX_DATA_54_const_net_21;
wire   [7:0]     TX_DATA_55_const_net_21;
wire   [7:0]     TX_DATA_56_const_net_21;
wire   [7:0]     TX_DATA_57_const_net_21;
wire   [7:0]     TX_DATA_58_const_net_21;
wire   [7:0]     TX_DATA_59_const_net_21;
wire   [7:0]     TX_DATA_60_const_net_21;
wire   [7:0]     TX_DATA_61_const_net_21;
wire   [7:0]     TX_DATA_62_const_net_21;
wire   [7:0]     TX_DATA_63_const_net_21;
wire   [7:0]     TX_DATA_64_const_net_21;
wire   [7:0]     TX_DATA_65_const_net_21;
wire   [7:0]     TX_DATA_66_const_net_21;
wire   [7:0]     TX_DATA_67_const_net_21;
wire   [7:0]     TX_DATA_68_const_net_21;
wire   [7:0]     TX_DATA_69_const_net_21;
wire   [7:0]     TX_DATA_70_const_net_21;
wire   [7:0]     TX_DATA_71_const_net_21;
wire   [7:0]     TX_DATA_72_const_net_21;
wire   [7:0]     TX_DATA_73_const_net_21;
wire   [7:0]     TX_DATA_74_const_net_21;
wire   [7:0]     TX_DATA_75_const_net_21;
wire   [7:0]     TX_DATA_76_const_net_21;
wire   [7:0]     TX_DATA_77_const_net_21;
wire   [7:0]     TX_DATA_78_const_net_21;
wire   [7:0]     TX_DATA_79_const_net_21;
wire   [7:0]     TX_DATA_80_const_net_21;
wire   [7:0]     TX_DATA_81_const_net_21;
wire   [7:0]     TX_DATA_82_const_net_21;
wire   [7:0]     TX_DATA_83_const_net_21;
wire   [7:0]     TX_DATA_84_const_net_21;
wire   [7:0]     TX_DATA_85_const_net_21;
wire   [7:0]     TX_DATA_86_const_net_21;
wire   [7:0]     TX_DATA_87_const_net_21;
wire   [7:0]     TX_DATA_88_const_net_21;
wire   [7:0]     TX_DATA_89_const_net_21;
wire   [7:0]     TX_DATA_90_const_net_21;
wire   [7:0]     TX_DATA_91_const_net_21;
wire   [7:0]     TX_DATA_92_const_net_21;
wire   [7:0]     TX_DATA_93_const_net_21;
wire   [7:0]     TX_DATA_94_const_net_21;
wire   [7:0]     TX_DATA_95_const_net_21;
wire   [7:0]     TX_DATA_96_const_net_21;
wire   [7:0]     TX_DATA_97_const_net_21;
wire   [7:0]     TX_DATA_98_const_net_21;
wire   [7:0]     TX_DATA_99_const_net_21;
wire   [7:0]     TX_DATA_100_const_net_21;
wire   [7:0]     TX_DATA_101_const_net_21;
wire   [7:0]     TX_DATA_102_const_net_21;
wire   [7:0]     TX_DATA_103_const_net_21;
wire   [7:0]     TX_DATA_104_const_net_21;
wire   [7:0]     TX_DATA_105_const_net_21;
wire   [7:0]     TX_DATA_106_const_net_21;
wire   [7:0]     TX_DATA_107_const_net_21;
wire   [7:0]     TX_DATA_108_const_net_21;
wire   [7:0]     TX_DATA_109_const_net_21;
wire   [7:0]     TX_DATA_110_const_net_21;
wire   [7:0]     TX_DATA_111_const_net_21;
wire   [7:0]     TX_DATA_112_const_net_21;
wire   [7:0]     TX_DATA_113_const_net_21;
wire   [7:0]     TX_DATA_114_const_net_21;
wire   [7:0]     TX_DATA_115_const_net_21;
wire   [7:0]     TX_DATA_116_const_net_21;
wire   [7:0]     TX_DATA_117_const_net_21;
wire   [7:0]     TX_DATA_118_const_net_21;
wire   [7:0]     TX_DATA_119_const_net_21;
wire   [7:0]     TX_DATA_120_const_net_21;
wire   [7:0]     TX_DATA_121_const_net_21;
wire   [7:0]     TX_DATA_122_const_net_21;
wire   [7:0]     TX_DATA_123_const_net_21;
wire   [7:0]     TX_DATA_124_const_net_21;
wire   [7:0]     TX_DATA_125_const_net_21;
wire   [7:0]     TX_DATA_126_const_net_21;
wire   [7:0]     TX_DATA_127_const_net_21;
wire   [3:0]     OE_DATA_8_const_net_21;
wire   [3:0]     OE_DATA_9_const_net_21;
wire   [3:0]     OE_DATA_10_const_net_21;
wire   [3:0]     OE_DATA_11_const_net_21;
wire   [3:0]     OE_DATA_12_const_net_21;
wire   [3:0]     OE_DATA_13_const_net_21;
wire   [3:0]     OE_DATA_14_const_net_21;
wire   [3:0]     OE_DATA_15_const_net_21;
wire   [3:0]     OE_DATA_16_const_net_21;
wire   [3:0]     OE_DATA_17_const_net_21;
wire   [3:0]     OE_DATA_18_const_net_21;
wire   [3:0]     OE_DATA_19_const_net_21;
wire   [3:0]     OE_DATA_20_const_net_21;
wire   [3:0]     OE_DATA_21_const_net_21;
wire   [3:0]     OE_DATA_22_const_net_21;
wire   [3:0]     OE_DATA_23_const_net_21;
wire   [3:0]     OE_DATA_24_const_net_21;
wire   [3:0]     OE_DATA_25_const_net_21;
wire   [3:0]     OE_DATA_26_const_net_21;
wire   [3:0]     OE_DATA_27_const_net_21;
wire   [3:0]     OE_DATA_28_const_net_21;
wire   [3:0]     OE_DATA_29_const_net_21;
wire   [3:0]     OE_DATA_30_const_net_21;
wire   [3:0]     OE_DATA_31_const_net_21;
wire   [3:0]     OE_DATA_32_const_net_21;
wire   [3:0]     OE_DATA_33_const_net_21;
wire   [3:0]     OE_DATA_34_const_net_21;
wire   [3:0]     OE_DATA_35_const_net_21;
wire   [3:0]     OE_DATA_36_const_net_21;
wire   [3:0]     OE_DATA_37_const_net_21;
wire   [3:0]     OE_DATA_38_const_net_21;
wire   [3:0]     OE_DATA_39_const_net_21;
wire   [3:0]     OE_DATA_40_const_net_21;
wire   [3:0]     OE_DATA_41_const_net_21;
wire   [3:0]     OE_DATA_42_const_net_21;
wire   [3:0]     OE_DATA_43_const_net_21;
wire   [3:0]     OE_DATA_44_const_net_21;
wire   [3:0]     OE_DATA_45_const_net_21;
wire   [3:0]     OE_DATA_46_const_net_21;
wire   [3:0]     OE_DATA_47_const_net_21;
wire   [3:0]     OE_DATA_48_const_net_21;
wire   [3:0]     OE_DATA_49_const_net_21;
wire   [3:0]     OE_DATA_50_const_net_21;
wire   [3:0]     OE_DATA_51_const_net_21;
wire   [3:0]     OE_DATA_52_const_net_21;
wire   [3:0]     OE_DATA_53_const_net_21;
wire   [3:0]     OE_DATA_54_const_net_21;
wire   [3:0]     OE_DATA_55_const_net_21;
wire   [3:0]     OE_DATA_56_const_net_21;
wire   [3:0]     OE_DATA_57_const_net_21;
wire   [3:0]     OE_DATA_58_const_net_21;
wire   [3:0]     OE_DATA_59_const_net_21;
wire   [3:0]     OE_DATA_60_const_net_21;
wire   [3:0]     OE_DATA_61_const_net_21;
wire   [3:0]     OE_DATA_62_const_net_21;
wire   [3:0]     OE_DATA_63_const_net_21;
wire   [3:0]     OE_DATA_64_const_net_21;
wire   [3:0]     OE_DATA_65_const_net_21;
wire   [3:0]     OE_DATA_66_const_net_21;
wire   [3:0]     OE_DATA_67_const_net_21;
wire   [3:0]     OE_DATA_68_const_net_21;
wire   [3:0]     OE_DATA_69_const_net_21;
wire   [3:0]     OE_DATA_70_const_net_21;
wire   [3:0]     OE_DATA_71_const_net_21;
wire   [3:0]     OE_DATA_72_const_net_21;
wire   [3:0]     OE_DATA_73_const_net_21;
wire   [3:0]     OE_DATA_74_const_net_21;
wire   [3:0]     OE_DATA_75_const_net_21;
wire   [3:0]     OE_DATA_76_const_net_21;
wire   [3:0]     OE_DATA_77_const_net_21;
wire   [3:0]     OE_DATA_78_const_net_21;
wire   [3:0]     OE_DATA_79_const_net_21;
wire   [3:0]     OE_DATA_80_const_net_21;
wire   [3:0]     OE_DATA_81_const_net_21;
wire   [3:0]     OE_DATA_82_const_net_21;
wire   [3:0]     OE_DATA_83_const_net_21;
wire   [3:0]     OE_DATA_84_const_net_21;
wire   [3:0]     OE_DATA_85_const_net_21;
wire   [3:0]     OE_DATA_86_const_net_21;
wire   [3:0]     OE_DATA_87_const_net_21;
wire   [3:0]     OE_DATA_88_const_net_21;
wire   [3:0]     OE_DATA_89_const_net_21;
wire   [3:0]     OE_DATA_90_const_net_21;
wire   [3:0]     OE_DATA_91_const_net_21;
wire   [3:0]     OE_DATA_92_const_net_21;
wire   [3:0]     OE_DATA_93_const_net_21;
wire   [3:0]     OE_DATA_94_const_net_21;
wire   [3:0]     OE_DATA_95_const_net_21;
wire   [3:0]     OE_DATA_96_const_net_21;
wire   [3:0]     OE_DATA_97_const_net_21;
wire   [3:0]     OE_DATA_98_const_net_21;
wire   [3:0]     OE_DATA_99_const_net_21;
wire   [3:0]     OE_DATA_100_const_net_21;
wire   [3:0]     OE_DATA_101_const_net_21;
wire   [3:0]     OE_DATA_102_const_net_21;
wire   [3:0]     OE_DATA_103_const_net_21;
wire   [3:0]     OE_DATA_104_const_net_21;
wire   [3:0]     OE_DATA_105_const_net_21;
wire   [3:0]     OE_DATA_106_const_net_21;
wire   [3:0]     OE_DATA_107_const_net_21;
wire   [3:0]     OE_DATA_108_const_net_21;
wire   [3:0]     OE_DATA_109_const_net_21;
wire   [3:0]     OE_DATA_110_const_net_21;
wire   [3:0]     OE_DATA_111_const_net_21;
wire   [3:0]     OE_DATA_112_const_net_21;
wire   [3:0]     OE_DATA_113_const_net_21;
wire   [3:0]     OE_DATA_114_const_net_21;
wire   [3:0]     OE_DATA_115_const_net_21;
wire   [3:0]     OE_DATA_116_const_net_21;
wire   [3:0]     OE_DATA_117_const_net_21;
wire   [3:0]     OE_DATA_118_const_net_21;
wire   [3:0]     OE_DATA_119_const_net_21;
wire   [3:0]     OE_DATA_120_const_net_21;
wire   [3:0]     OE_DATA_121_const_net_21;
wire   [3:0]     OE_DATA_122_const_net_21;
wire   [3:0]     OE_DATA_123_const_net_21;
wire   [3:0]     OE_DATA_124_const_net_21;
wire   [3:0]     OE_DATA_125_const_net_21;
wire   [3:0]     OE_DATA_126_const_net_21;
wire   [3:0]     OE_DATA_127_const_net_21;
wire   [7:0]     PAD_I_const_net_4;
wire   [7:0]     PAD_N_const_net_4;
wire   [7:0]     PAD_I_N_const_net_4;
wire   [7:0]     TX_DATA_1_const_net_17;
wire   [7:0]     TX_DATA_2_const_net_19;
wire   [7:0]     TX_DATA_3_const_net_19;
wire   [7:0]     TX_DATA_4_const_net_19;
wire   [7:0]     TX_DATA_5_const_net_19;
wire   [7:0]     TX_DATA_6_const_net_19;
wire   [7:0]     TX_DATA_7_const_net_19;
wire   [7:0]     TX_DATA_8_const_net_21;
wire   [7:0]     TX_DATA_9_const_net_21;
wire   [7:0]     TX_DATA_10_const_net_21;
wire   [7:0]     TX_DATA_11_const_net_21;
wire   [7:0]     TX_DATA_12_const_net_22;
wire   [7:0]     TX_DATA_13_const_net_22;
wire   [7:0]     TX_DATA_14_const_net_22;
wire   [7:0]     TX_DATA_15_const_net_22;
wire   [7:0]     TX_DATA_16_const_net_22;
wire   [7:0]     TX_DATA_17_const_net_22;
wire   [7:0]     TX_DATA_18_const_net_22;
wire   [7:0]     TX_DATA_19_const_net_22;
wire   [7:0]     TX_DATA_20_const_net_22;
wire   [7:0]     TX_DATA_21_const_net_22;
wire   [7:0]     TX_DATA_22_const_net_22;
wire   [7:0]     TX_DATA_23_const_net_22;
wire   [7:0]     TX_DATA_24_const_net_22;
wire   [7:0]     TX_DATA_25_const_net_22;
wire   [7:0]     TX_DATA_26_const_net_22;
wire   [7:0]     TX_DATA_27_const_net_22;
wire   [7:0]     TX_DATA_28_const_net_22;
wire   [7:0]     TX_DATA_29_const_net_22;
wire   [7:0]     TX_DATA_30_const_net_22;
wire   [7:0]     TX_DATA_31_const_net_22;
wire   [7:0]     TX_DATA_32_const_net_22;
wire   [7:0]     TX_DATA_33_const_net_22;
wire   [7:0]     TX_DATA_34_const_net_22;
wire   [7:0]     TX_DATA_35_const_net_22;
wire   [7:0]     TX_DATA_36_const_net_22;
wire   [7:0]     TX_DATA_37_const_net_22;
wire   [7:0]     TX_DATA_38_const_net_22;
wire   [7:0]     TX_DATA_39_const_net_22;
wire   [7:0]     TX_DATA_40_const_net_22;
wire   [7:0]     TX_DATA_41_const_net_22;
wire   [7:0]     TX_DATA_42_const_net_22;
wire   [7:0]     TX_DATA_43_const_net_22;
wire   [7:0]     TX_DATA_44_const_net_22;
wire   [7:0]     TX_DATA_45_const_net_22;
wire   [7:0]     TX_DATA_46_const_net_22;
wire   [7:0]     TX_DATA_47_const_net_22;
wire   [7:0]     TX_DATA_48_const_net_22;
wire   [7:0]     TX_DATA_49_const_net_22;
wire   [7:0]     TX_DATA_50_const_net_22;
wire   [7:0]     TX_DATA_51_const_net_22;
wire   [7:0]     TX_DATA_52_const_net_22;
wire   [7:0]     TX_DATA_53_const_net_22;
wire   [7:0]     TX_DATA_54_const_net_22;
wire   [7:0]     TX_DATA_55_const_net_22;
wire   [7:0]     TX_DATA_56_const_net_22;
wire   [7:0]     TX_DATA_57_const_net_22;
wire   [7:0]     TX_DATA_58_const_net_22;
wire   [7:0]     TX_DATA_59_const_net_22;
wire   [7:0]     TX_DATA_60_const_net_22;
wire   [7:0]     TX_DATA_61_const_net_22;
wire   [7:0]     TX_DATA_62_const_net_22;
wire   [7:0]     TX_DATA_63_const_net_22;
wire   [7:0]     TX_DATA_64_const_net_22;
wire   [7:0]     TX_DATA_65_const_net_22;
wire   [7:0]     TX_DATA_66_const_net_22;
wire   [7:0]     TX_DATA_67_const_net_22;
wire   [7:0]     TX_DATA_68_const_net_22;
wire   [7:0]     TX_DATA_69_const_net_22;
wire   [7:0]     TX_DATA_70_const_net_22;
wire   [7:0]     TX_DATA_71_const_net_22;
wire   [7:0]     TX_DATA_72_const_net_22;
wire   [7:0]     TX_DATA_73_const_net_22;
wire   [7:0]     TX_DATA_74_const_net_22;
wire   [7:0]     TX_DATA_75_const_net_22;
wire   [7:0]     TX_DATA_76_const_net_22;
wire   [7:0]     TX_DATA_77_const_net_22;
wire   [7:0]     TX_DATA_78_const_net_22;
wire   [7:0]     TX_DATA_79_const_net_22;
wire   [7:0]     TX_DATA_80_const_net_22;
wire   [7:0]     TX_DATA_81_const_net_22;
wire   [7:0]     TX_DATA_82_const_net_22;
wire   [7:0]     TX_DATA_83_const_net_22;
wire   [7:0]     TX_DATA_84_const_net_22;
wire   [7:0]     TX_DATA_85_const_net_22;
wire   [7:0]     TX_DATA_86_const_net_22;
wire   [7:0]     TX_DATA_87_const_net_22;
wire   [7:0]     TX_DATA_88_const_net_22;
wire   [7:0]     TX_DATA_89_const_net_22;
wire   [7:0]     TX_DATA_90_const_net_22;
wire   [7:0]     TX_DATA_91_const_net_22;
wire   [7:0]     TX_DATA_92_const_net_22;
wire   [7:0]     TX_DATA_93_const_net_22;
wire   [7:0]     TX_DATA_94_const_net_22;
wire   [7:0]     TX_DATA_95_const_net_22;
wire   [7:0]     TX_DATA_96_const_net_22;
wire   [7:0]     TX_DATA_97_const_net_22;
wire   [7:0]     TX_DATA_98_const_net_22;
wire   [7:0]     TX_DATA_99_const_net_22;
wire   [7:0]     TX_DATA_100_const_net_22;
wire   [7:0]     TX_DATA_101_const_net_22;
wire   [7:0]     TX_DATA_102_const_net_22;
wire   [7:0]     TX_DATA_103_const_net_22;
wire   [7:0]     TX_DATA_104_const_net_22;
wire   [7:0]     TX_DATA_105_const_net_22;
wire   [7:0]     TX_DATA_106_const_net_22;
wire   [7:0]     TX_DATA_107_const_net_22;
wire   [7:0]     TX_DATA_108_const_net_22;
wire   [7:0]     TX_DATA_109_const_net_22;
wire   [7:0]     TX_DATA_110_const_net_22;
wire   [7:0]     TX_DATA_111_const_net_22;
wire   [7:0]     TX_DATA_112_const_net_22;
wire   [7:0]     TX_DATA_113_const_net_22;
wire   [7:0]     TX_DATA_114_const_net_22;
wire   [7:0]     TX_DATA_115_const_net_22;
wire   [7:0]     TX_DATA_116_const_net_22;
wire   [7:0]     TX_DATA_117_const_net_22;
wire   [7:0]     TX_DATA_118_const_net_22;
wire   [7:0]     TX_DATA_119_const_net_22;
wire   [7:0]     TX_DATA_120_const_net_22;
wire   [7:0]     TX_DATA_121_const_net_22;
wire   [7:0]     TX_DATA_122_const_net_22;
wire   [7:0]     TX_DATA_123_const_net_22;
wire   [7:0]     TX_DATA_124_const_net_22;
wire   [7:0]     TX_DATA_125_const_net_22;
wire   [7:0]     TX_DATA_126_const_net_22;
wire   [7:0]     TX_DATA_127_const_net_22;
wire   [3:0]     OE_DATA_1_const_net_20;
wire   [3:0]     OE_DATA_2_const_net_20;
wire   [3:0]     OE_DATA_3_const_net_20;
wire   [3:0]     OE_DATA_4_const_net_20;
wire   [3:0]     OE_DATA_5_const_net_20;
wire   [3:0]     OE_DATA_6_const_net_20;
wire   [3:0]     OE_DATA_7_const_net_20;
wire   [3:0]     OE_DATA_8_const_net_22;
wire   [3:0]     OE_DATA_9_const_net_22;
wire   [3:0]     OE_DATA_10_const_net_22;
wire   [3:0]     OE_DATA_11_const_net_22;
wire   [3:0]     OE_DATA_12_const_net_22;
wire   [3:0]     OE_DATA_13_const_net_22;
wire   [3:0]     OE_DATA_14_const_net_22;
wire   [3:0]     OE_DATA_15_const_net_22;
wire   [3:0]     OE_DATA_16_const_net_22;
wire   [3:0]     OE_DATA_17_const_net_22;
wire   [3:0]     OE_DATA_18_const_net_22;
wire   [3:0]     OE_DATA_19_const_net_22;
wire   [3:0]     OE_DATA_20_const_net_22;
wire   [3:0]     OE_DATA_21_const_net_22;
wire   [3:0]     OE_DATA_22_const_net_22;
wire   [3:0]     OE_DATA_23_const_net_22;
wire   [3:0]     OE_DATA_24_const_net_22;
wire   [3:0]     OE_DATA_25_const_net_22;
wire   [3:0]     OE_DATA_26_const_net_22;
wire   [3:0]     OE_DATA_27_const_net_22;
wire   [3:0]     OE_DATA_28_const_net_22;
wire   [3:0]     OE_DATA_29_const_net_22;
wire   [3:0]     OE_DATA_30_const_net_22;
wire   [3:0]     OE_DATA_31_const_net_22;
wire   [3:0]     OE_DATA_32_const_net_22;
wire   [3:0]     OE_DATA_33_const_net_22;
wire   [3:0]     OE_DATA_34_const_net_22;
wire   [3:0]     OE_DATA_35_const_net_22;
wire   [3:0]     OE_DATA_36_const_net_22;
wire   [3:0]     OE_DATA_37_const_net_22;
wire   [3:0]     OE_DATA_38_const_net_22;
wire   [3:0]     OE_DATA_39_const_net_22;
wire   [3:0]     OE_DATA_40_const_net_22;
wire   [3:0]     OE_DATA_41_const_net_22;
wire   [3:0]     OE_DATA_42_const_net_22;
wire   [3:0]     OE_DATA_43_const_net_22;
wire   [3:0]     OE_DATA_44_const_net_22;
wire   [3:0]     OE_DATA_45_const_net_22;
wire   [3:0]     OE_DATA_46_const_net_22;
wire   [3:0]     OE_DATA_47_const_net_22;
wire   [3:0]     OE_DATA_48_const_net_22;
wire   [3:0]     OE_DATA_49_const_net_22;
wire   [3:0]     OE_DATA_50_const_net_22;
wire   [3:0]     OE_DATA_51_const_net_22;
wire   [3:0]     OE_DATA_52_const_net_22;
wire   [3:0]     OE_DATA_53_const_net_22;
wire   [3:0]     OE_DATA_54_const_net_22;
wire   [3:0]     OE_DATA_55_const_net_22;
wire   [3:0]     OE_DATA_56_const_net_22;
wire   [3:0]     OE_DATA_57_const_net_22;
wire   [3:0]     OE_DATA_58_const_net_22;
wire   [3:0]     OE_DATA_59_const_net_22;
wire   [3:0]     OE_DATA_60_const_net_22;
wire   [3:0]     OE_DATA_61_const_net_22;
wire   [3:0]     OE_DATA_62_const_net_22;
wire   [3:0]     OE_DATA_63_const_net_22;
wire   [3:0]     OE_DATA_64_const_net_22;
wire   [3:0]     OE_DATA_65_const_net_22;
wire   [3:0]     OE_DATA_66_const_net_22;
wire   [3:0]     OE_DATA_67_const_net_22;
wire   [3:0]     OE_DATA_68_const_net_22;
wire   [3:0]     OE_DATA_69_const_net_22;
wire   [3:0]     OE_DATA_70_const_net_22;
wire   [3:0]     OE_DATA_71_const_net_22;
wire   [3:0]     OE_DATA_72_const_net_22;
wire   [3:0]     OE_DATA_73_const_net_22;
wire   [3:0]     OE_DATA_74_const_net_22;
wire   [3:0]     OE_DATA_75_const_net_22;
wire   [3:0]     OE_DATA_76_const_net_22;
wire   [3:0]     OE_DATA_77_const_net_22;
wire   [3:0]     OE_DATA_78_const_net_22;
wire   [3:0]     OE_DATA_79_const_net_22;
wire   [3:0]     OE_DATA_80_const_net_22;
wire   [3:0]     OE_DATA_81_const_net_22;
wire   [3:0]     OE_DATA_82_const_net_22;
wire   [3:0]     OE_DATA_83_const_net_22;
wire   [3:0]     OE_DATA_84_const_net_22;
wire   [3:0]     OE_DATA_85_const_net_22;
wire   [3:0]     OE_DATA_86_const_net_22;
wire   [3:0]     OE_DATA_87_const_net_22;
wire   [3:0]     OE_DATA_88_const_net_22;
wire   [3:0]     OE_DATA_89_const_net_22;
wire   [3:0]     OE_DATA_90_const_net_22;
wire   [3:0]     OE_DATA_91_const_net_22;
wire   [3:0]     OE_DATA_92_const_net_22;
wire   [3:0]     OE_DATA_93_const_net_22;
wire   [3:0]     OE_DATA_94_const_net_22;
wire   [3:0]     OE_DATA_95_const_net_22;
wire   [3:0]     OE_DATA_96_const_net_22;
wire   [3:0]     OE_DATA_97_const_net_22;
wire   [3:0]     OE_DATA_98_const_net_22;
wire   [3:0]     OE_DATA_99_const_net_22;
wire   [3:0]     OE_DATA_100_const_net_22;
wire   [3:0]     OE_DATA_101_const_net_22;
wire   [3:0]     OE_DATA_102_const_net_22;
wire   [3:0]     OE_DATA_103_const_net_22;
wire   [3:0]     OE_DATA_104_const_net_22;
wire   [3:0]     OE_DATA_105_const_net_22;
wire   [3:0]     OE_DATA_106_const_net_22;
wire   [3:0]     OE_DATA_107_const_net_22;
wire   [3:0]     OE_DATA_108_const_net_22;
wire   [3:0]     OE_DATA_109_const_net_22;
wire   [3:0]     OE_DATA_110_const_net_22;
wire   [3:0]     OE_DATA_111_const_net_22;
wire   [3:0]     OE_DATA_112_const_net_22;
wire   [3:0]     OE_DATA_113_const_net_22;
wire   [3:0]     OE_DATA_114_const_net_22;
wire   [3:0]     OE_DATA_115_const_net_22;
wire   [3:0]     OE_DATA_116_const_net_22;
wire   [3:0]     OE_DATA_117_const_net_22;
wire   [3:0]     OE_DATA_118_const_net_22;
wire   [3:0]     OE_DATA_119_const_net_22;
wire   [3:0]     OE_DATA_120_const_net_22;
wire   [3:0]     OE_DATA_121_const_net_22;
wire   [3:0]     OE_DATA_122_const_net_22;
wire   [3:0]     OE_DATA_123_const_net_22;
wire   [3:0]     OE_DATA_124_const_net_22;
wire   [3:0]     OE_DATA_125_const_net_22;
wire   [3:0]     OE_DATA_126_const_net_22;
wire   [3:0]     OE_DATA_127_const_net_22;
wire   [1:0]     RX_DQS_90_const_net_17;
wire   [2:0]     FIFO_WR_PTR_const_net_18;
wire   [2:0]     FIFO_RD_PTR_const_net_18;
wire   [2:0]     EYE_MONITOR_LANE_WIDTH_const_net_19;
wire   [1:0]     TX_DATA_1_const_net_18;
wire   [1:0]     TX_DATA_2_const_net_20;
wire   [1:0]     TX_DATA_3_const_net_20;
wire   [1:0]     TX_DATA_4_const_net_20;
wire   [1:0]     TX_DATA_5_const_net_20;
wire   [1:0]     TX_DATA_6_const_net_20;
wire   [1:0]     TX_DATA_7_const_net_20;
wire   [1:0]     TX_DATA_8_const_net_22;
wire   [1:0]     TX_DATA_9_const_net_22;
wire   [1:0]     TX_DATA_10_const_net_22;
wire   [1:0]     TX_DATA_11_const_net_22;
wire   [1:0]     TX_DATA_12_const_net_23;
wire   [1:0]     TX_DATA_13_const_net_23;
wire   [1:0]     TX_DATA_14_const_net_23;
wire   [1:0]     TX_DATA_15_const_net_23;
wire   [1:0]     TX_DATA_16_const_net_23;
wire   [1:0]     TX_DATA_17_const_net_23;
wire   [1:0]     TX_DATA_18_const_net_23;
wire   [1:0]     TX_DATA_19_const_net_23;
wire   [1:0]     TX_DATA_20_const_net_23;
wire   [1:0]     TX_DATA_21_const_net_23;
wire   [1:0]     TX_DATA_22_const_net_23;
wire   [1:0]     TX_DATA_23_const_net_23;
wire   [1:0]     TX_DATA_24_const_net_23;
wire   [1:0]     TX_DATA_25_const_net_23;
wire   [1:0]     TX_DATA_26_const_net_23;
wire   [1:0]     TX_DATA_27_const_net_23;
wire   [1:0]     TX_DATA_28_const_net_23;
wire   [1:0]     TX_DATA_29_const_net_23;
wire   [1:0]     TX_DATA_30_const_net_23;
wire   [1:0]     TX_DATA_31_const_net_23;
wire   [1:0]     TX_DATA_32_const_net_23;
wire   [1:0]     TX_DATA_33_const_net_23;
wire   [1:0]     TX_DATA_34_const_net_23;
wire   [1:0]     TX_DATA_35_const_net_23;
wire   [1:0]     TX_DATA_36_const_net_23;
wire   [1:0]     TX_DATA_37_const_net_23;
wire   [1:0]     TX_DATA_38_const_net_23;
wire   [1:0]     TX_DATA_39_const_net_23;
wire   [1:0]     TX_DATA_40_const_net_23;
wire   [1:0]     TX_DATA_41_const_net_23;
wire   [1:0]     TX_DATA_42_const_net_23;
wire   [1:0]     TX_DATA_43_const_net_23;
wire   [1:0]     TX_DATA_44_const_net_23;
wire   [1:0]     TX_DATA_45_const_net_23;
wire   [1:0]     TX_DATA_46_const_net_23;
wire   [1:0]     TX_DATA_47_const_net_23;
wire   [1:0]     TX_DATA_48_const_net_23;
wire   [1:0]     TX_DATA_49_const_net_23;
wire   [1:0]     TX_DATA_50_const_net_23;
wire   [1:0]     TX_DATA_51_const_net_23;
wire   [1:0]     TX_DATA_52_const_net_23;
wire   [1:0]     TX_DATA_53_const_net_23;
wire   [1:0]     TX_DATA_54_const_net_23;
wire   [1:0]     TX_DATA_55_const_net_23;
wire   [1:0]     TX_DATA_56_const_net_23;
wire   [1:0]     TX_DATA_57_const_net_23;
wire   [1:0]     TX_DATA_58_const_net_23;
wire   [1:0]     TX_DATA_59_const_net_23;
wire   [1:0]     TX_DATA_60_const_net_23;
wire   [1:0]     TX_DATA_61_const_net_23;
wire   [1:0]     TX_DATA_62_const_net_23;
wire   [1:0]     TX_DATA_63_const_net_23;
wire   [1:0]     TX_DATA_64_const_net_23;
wire   [1:0]     TX_DATA_65_const_net_23;
wire   [1:0]     TX_DATA_66_const_net_23;
wire   [1:0]     TX_DATA_67_const_net_23;
wire   [1:0]     TX_DATA_68_const_net_23;
wire   [1:0]     TX_DATA_69_const_net_23;
wire   [1:0]     TX_DATA_70_const_net_23;
wire   [1:0]     TX_DATA_71_const_net_23;
wire   [1:0]     TX_DATA_72_const_net_23;
wire   [1:0]     TX_DATA_73_const_net_23;
wire   [1:0]     TX_DATA_74_const_net_23;
wire   [1:0]     TX_DATA_75_const_net_23;
wire   [1:0]     TX_DATA_76_const_net_23;
wire   [1:0]     TX_DATA_77_const_net_23;
wire   [1:0]     TX_DATA_78_const_net_23;
wire   [1:0]     TX_DATA_79_const_net_23;
wire   [1:0]     TX_DATA_80_const_net_23;
wire   [1:0]     TX_DATA_81_const_net_23;
wire   [1:0]     TX_DATA_82_const_net_23;
wire   [1:0]     TX_DATA_83_const_net_23;
wire   [1:0]     TX_DATA_84_const_net_23;
wire   [1:0]     TX_DATA_85_const_net_23;
wire   [1:0]     TX_DATA_86_const_net_23;
wire   [1:0]     TX_DATA_87_const_net_23;
wire   [1:0]     TX_DATA_88_const_net_23;
wire   [1:0]     TX_DATA_89_const_net_23;
wire   [1:0]     TX_DATA_90_const_net_23;
wire   [1:0]     TX_DATA_91_const_net_23;
wire   [1:0]     TX_DATA_92_const_net_23;
wire   [1:0]     TX_DATA_93_const_net_23;
wire   [1:0]     TX_DATA_94_const_net_23;
wire   [1:0]     TX_DATA_95_const_net_23;
wire   [1:0]     TX_DATA_96_const_net_23;
wire   [1:0]     TX_DATA_97_const_net_23;
wire   [1:0]     TX_DATA_98_const_net_23;
wire   [1:0]     TX_DATA_99_const_net_23;
wire   [1:0]     TX_DATA_100_const_net_23;
wire   [1:0]     TX_DATA_101_const_net_23;
wire   [1:0]     TX_DATA_102_const_net_23;
wire   [1:0]     TX_DATA_103_const_net_23;
wire   [1:0]     TX_DATA_104_const_net_23;
wire   [1:0]     TX_DATA_105_const_net_23;
wire   [1:0]     TX_DATA_106_const_net_23;
wire   [1:0]     TX_DATA_107_const_net_23;
wire   [1:0]     TX_DATA_108_const_net_23;
wire   [1:0]     TX_DATA_109_const_net_23;
wire   [1:0]     TX_DATA_110_const_net_23;
wire   [1:0]     TX_DATA_111_const_net_23;
wire   [1:0]     TX_DATA_112_const_net_23;
wire   [1:0]     TX_DATA_113_const_net_23;
wire   [1:0]     TX_DATA_114_const_net_23;
wire   [1:0]     TX_DATA_115_const_net_23;
wire   [1:0]     TX_DATA_116_const_net_23;
wire   [1:0]     TX_DATA_117_const_net_23;
wire   [1:0]     TX_DATA_118_const_net_23;
wire   [1:0]     TX_DATA_119_const_net_23;
wire   [1:0]     TX_DATA_120_const_net_23;
wire   [1:0]     TX_DATA_121_const_net_23;
wire   [1:0]     TX_DATA_122_const_net_23;
wire   [1:0]     TX_DATA_123_const_net_23;
wire   [1:0]     TX_DATA_124_const_net_23;
wire   [1:0]     TX_DATA_125_const_net_23;
wire   [1:0]     TX_DATA_126_const_net_23;
wire   [1:0]     TX_DATA_127_const_net_23;
wire   [1:0]     OE_DATA_1_const_net_21;
wire   [1:0]     OE_DATA_2_const_net_21;
wire   [1:0]     OE_DATA_3_const_net_21;
wire   [1:0]     OE_DATA_4_const_net_21;
wire   [1:0]     OE_DATA_5_const_net_21;
wire   [1:0]     OE_DATA_6_const_net_21;
wire   [1:0]     OE_DATA_7_const_net_21;
wire   [1:0]     OE_DATA_8_const_net_23;
wire   [1:0]     OE_DATA_9_const_net_23;
wire   [1:0]     OE_DATA_10_const_net_23;
wire   [1:0]     OE_DATA_11_const_net_23;
wire   [1:0]     OE_DATA_12_const_net_23;
wire   [1:0]     OE_DATA_13_const_net_23;
wire   [1:0]     OE_DATA_14_const_net_23;
wire   [1:0]     OE_DATA_15_const_net_23;
wire   [1:0]     OE_DATA_16_const_net_23;
wire   [1:0]     OE_DATA_17_const_net_23;
wire   [1:0]     OE_DATA_18_const_net_23;
wire   [1:0]     OE_DATA_19_const_net_23;
wire   [1:0]     OE_DATA_20_const_net_23;
wire   [1:0]     OE_DATA_21_const_net_23;
wire   [1:0]     OE_DATA_22_const_net_23;
wire   [1:0]     OE_DATA_23_const_net_23;
wire   [1:0]     OE_DATA_24_const_net_23;
wire   [1:0]     OE_DATA_25_const_net_23;
wire   [1:0]     OE_DATA_26_const_net_23;
wire   [1:0]     OE_DATA_27_const_net_23;
wire   [1:0]     OE_DATA_28_const_net_23;
wire   [1:0]     OE_DATA_29_const_net_23;
wire   [1:0]     OE_DATA_30_const_net_23;
wire   [1:0]     OE_DATA_31_const_net_23;
wire   [1:0]     OE_DATA_32_const_net_23;
wire   [1:0]     OE_DATA_33_const_net_23;
wire   [1:0]     OE_DATA_34_const_net_23;
wire   [1:0]     OE_DATA_35_const_net_23;
wire   [1:0]     OE_DATA_36_const_net_23;
wire   [1:0]     OE_DATA_37_const_net_23;
wire   [1:0]     OE_DATA_38_const_net_23;
wire   [1:0]     OE_DATA_39_const_net_23;
wire   [1:0]     OE_DATA_40_const_net_23;
wire   [1:0]     OE_DATA_41_const_net_23;
wire   [1:0]     OE_DATA_42_const_net_23;
wire   [1:0]     OE_DATA_43_const_net_23;
wire   [1:0]     OE_DATA_44_const_net_23;
wire   [1:0]     OE_DATA_45_const_net_23;
wire   [1:0]     OE_DATA_46_const_net_23;
wire   [1:0]     OE_DATA_47_const_net_23;
wire   [1:0]     OE_DATA_48_const_net_23;
wire   [1:0]     OE_DATA_49_const_net_23;
wire   [1:0]     OE_DATA_50_const_net_23;
wire   [1:0]     OE_DATA_51_const_net_23;
wire   [1:0]     OE_DATA_52_const_net_23;
wire   [1:0]     OE_DATA_53_const_net_23;
wire   [1:0]     OE_DATA_54_const_net_23;
wire   [1:0]     OE_DATA_55_const_net_23;
wire   [1:0]     OE_DATA_56_const_net_23;
wire   [1:0]     OE_DATA_57_const_net_23;
wire   [1:0]     OE_DATA_58_const_net_23;
wire   [1:0]     OE_DATA_59_const_net_23;
wire   [1:0]     OE_DATA_60_const_net_23;
wire   [1:0]     OE_DATA_61_const_net_23;
wire   [1:0]     OE_DATA_62_const_net_23;
wire   [1:0]     OE_DATA_63_const_net_23;
wire   [1:0]     OE_DATA_64_const_net_23;
wire   [1:0]     OE_DATA_65_const_net_23;
wire   [1:0]     OE_DATA_66_const_net_23;
wire   [1:0]     OE_DATA_67_const_net_23;
wire   [1:0]     OE_DATA_68_const_net_23;
wire   [1:0]     OE_DATA_69_const_net_23;
wire   [1:0]     OE_DATA_70_const_net_23;
wire   [1:0]     OE_DATA_71_const_net_23;
wire   [1:0]     OE_DATA_72_const_net_23;
wire   [1:0]     OE_DATA_73_const_net_23;
wire   [1:0]     OE_DATA_74_const_net_23;
wire   [1:0]     OE_DATA_75_const_net_23;
wire   [1:0]     OE_DATA_76_const_net_23;
wire   [1:0]     OE_DATA_77_const_net_23;
wire   [1:0]     OE_DATA_78_const_net_23;
wire   [1:0]     OE_DATA_79_const_net_23;
wire   [1:0]     OE_DATA_80_const_net_23;
wire   [1:0]     OE_DATA_81_const_net_23;
wire   [1:0]     OE_DATA_82_const_net_23;
wire   [1:0]     OE_DATA_83_const_net_23;
wire   [1:0]     OE_DATA_84_const_net_23;
wire   [1:0]     OE_DATA_85_const_net_23;
wire   [1:0]     OE_DATA_86_const_net_23;
wire   [1:0]     OE_DATA_87_const_net_23;
wire   [1:0]     OE_DATA_88_const_net_23;
wire   [1:0]     OE_DATA_89_const_net_23;
wire   [1:0]     OE_DATA_90_const_net_23;
wire   [1:0]     OE_DATA_91_const_net_23;
wire   [1:0]     OE_DATA_92_const_net_23;
wire   [1:0]     OE_DATA_93_const_net_23;
wire   [1:0]     OE_DATA_94_const_net_23;
wire   [1:0]     OE_DATA_95_const_net_23;
wire   [1:0]     OE_DATA_96_const_net_23;
wire   [1:0]     OE_DATA_97_const_net_23;
wire   [1:0]     OE_DATA_98_const_net_23;
wire   [1:0]     OE_DATA_99_const_net_23;
wire   [1:0]     OE_DATA_100_const_net_23;
wire   [1:0]     OE_DATA_101_const_net_23;
wire   [1:0]     OE_DATA_102_const_net_23;
wire   [1:0]     OE_DATA_103_const_net_23;
wire   [1:0]     OE_DATA_104_const_net_23;
wire   [1:0]     OE_DATA_105_const_net_23;
wire   [1:0]     OE_DATA_106_const_net_23;
wire   [1:0]     OE_DATA_107_const_net_23;
wire   [1:0]     OE_DATA_108_const_net_23;
wire   [1:0]     OE_DATA_109_const_net_23;
wire   [1:0]     OE_DATA_110_const_net_23;
wire   [1:0]     OE_DATA_111_const_net_23;
wire   [1:0]     OE_DATA_112_const_net_23;
wire   [1:0]     OE_DATA_113_const_net_23;
wire   [1:0]     OE_DATA_114_const_net_23;
wire   [1:0]     OE_DATA_115_const_net_23;
wire   [1:0]     OE_DATA_116_const_net_23;
wire   [1:0]     OE_DATA_117_const_net_23;
wire   [1:0]     OE_DATA_118_const_net_23;
wire   [1:0]     OE_DATA_119_const_net_23;
wire   [1:0]     OE_DATA_120_const_net_23;
wire   [1:0]     OE_DATA_121_const_net_23;
wire   [1:0]     OE_DATA_122_const_net_23;
wire   [1:0]     OE_DATA_123_const_net_23;
wire   [1:0]     OE_DATA_124_const_net_23;
wire   [1:0]     OE_DATA_125_const_net_23;
wire   [1:0]     OE_DATA_126_const_net_23;
wire   [1:0]     OE_DATA_127_const_net_23;
wire   [1:0]     RX_DQS_90_const_net_18;
wire   [2:0]     EYE_MONITOR_LANE_WIDTH_const_net_20;
wire   [7:0]     TX_DATA_1_const_net_19;
wire   [7:0]     TX_DATA_2_const_net_21;
wire   [7:0]     TX_DATA_3_const_net_21;
wire   [7:0]     TX_DATA_4_const_net_21;
wire   [7:0]     TX_DATA_5_const_net_21;
wire   [7:0]     TX_DATA_6_const_net_21;
wire   [7:0]     TX_DATA_7_const_net_21;
wire   [7:0]     TX_DATA_8_const_net_23;
wire   [7:0]     TX_DATA_9_const_net_23;
wire   [7:0]     TX_DATA_10_const_net_23;
wire   [7:0]     TX_DATA_11_const_net_23;
wire   [7:0]     TX_DATA_12_const_net_24;
wire   [7:0]     TX_DATA_13_const_net_24;
wire   [7:0]     TX_DATA_14_const_net_24;
wire   [7:0]     TX_DATA_15_const_net_24;
wire   [7:0]     TX_DATA_16_const_net_24;
wire   [7:0]     TX_DATA_17_const_net_24;
wire   [7:0]     TX_DATA_18_const_net_24;
wire   [7:0]     TX_DATA_19_const_net_24;
wire   [7:0]     TX_DATA_20_const_net_24;
wire   [7:0]     TX_DATA_21_const_net_24;
wire   [7:0]     TX_DATA_22_const_net_24;
wire   [7:0]     TX_DATA_23_const_net_24;
wire   [7:0]     TX_DATA_24_const_net_24;
wire   [7:0]     TX_DATA_25_const_net_24;
wire   [7:0]     TX_DATA_26_const_net_24;
wire   [7:0]     TX_DATA_27_const_net_24;
wire   [7:0]     TX_DATA_28_const_net_24;
wire   [7:0]     TX_DATA_29_const_net_24;
wire   [7:0]     TX_DATA_30_const_net_24;
wire   [7:0]     TX_DATA_31_const_net_24;
wire   [7:0]     TX_DATA_32_const_net_24;
wire   [7:0]     TX_DATA_33_const_net_24;
wire   [7:0]     TX_DATA_34_const_net_24;
wire   [7:0]     TX_DATA_35_const_net_24;
wire   [7:0]     TX_DATA_36_const_net_24;
wire   [7:0]     TX_DATA_37_const_net_24;
wire   [7:0]     TX_DATA_38_const_net_24;
wire   [7:0]     TX_DATA_39_const_net_24;
wire   [7:0]     TX_DATA_40_const_net_24;
wire   [7:0]     TX_DATA_41_const_net_24;
wire   [7:0]     TX_DATA_42_const_net_24;
wire   [7:0]     TX_DATA_43_const_net_24;
wire   [7:0]     TX_DATA_44_const_net_24;
wire   [7:0]     TX_DATA_45_const_net_24;
wire   [7:0]     TX_DATA_46_const_net_24;
wire   [7:0]     TX_DATA_47_const_net_24;
wire   [7:0]     TX_DATA_48_const_net_24;
wire   [7:0]     TX_DATA_49_const_net_24;
wire   [7:0]     TX_DATA_50_const_net_24;
wire   [7:0]     TX_DATA_51_const_net_24;
wire   [7:0]     TX_DATA_52_const_net_24;
wire   [7:0]     TX_DATA_53_const_net_24;
wire   [7:0]     TX_DATA_54_const_net_24;
wire   [7:0]     TX_DATA_55_const_net_24;
wire   [7:0]     TX_DATA_56_const_net_24;
wire   [7:0]     TX_DATA_57_const_net_24;
wire   [7:0]     TX_DATA_58_const_net_24;
wire   [7:0]     TX_DATA_59_const_net_24;
wire   [7:0]     TX_DATA_60_const_net_24;
wire   [7:0]     TX_DATA_61_const_net_24;
wire   [7:0]     TX_DATA_62_const_net_24;
wire   [7:0]     TX_DATA_63_const_net_24;
wire   [7:0]     TX_DATA_64_const_net_24;
wire   [7:0]     TX_DATA_65_const_net_24;
wire   [7:0]     TX_DATA_66_const_net_24;
wire   [7:0]     TX_DATA_67_const_net_24;
wire   [7:0]     TX_DATA_68_const_net_24;
wire   [7:0]     TX_DATA_69_const_net_24;
wire   [7:0]     TX_DATA_70_const_net_24;
wire   [7:0]     TX_DATA_71_const_net_24;
wire   [7:0]     TX_DATA_72_const_net_24;
wire   [7:0]     TX_DATA_73_const_net_24;
wire   [7:0]     TX_DATA_74_const_net_24;
wire   [7:0]     TX_DATA_75_const_net_24;
wire   [7:0]     TX_DATA_76_const_net_24;
wire   [7:0]     TX_DATA_77_const_net_24;
wire   [7:0]     TX_DATA_78_const_net_24;
wire   [7:0]     TX_DATA_79_const_net_24;
wire   [7:0]     TX_DATA_80_const_net_24;
wire   [7:0]     TX_DATA_81_const_net_24;
wire   [7:0]     TX_DATA_82_const_net_24;
wire   [7:0]     TX_DATA_83_const_net_24;
wire   [7:0]     TX_DATA_84_const_net_24;
wire   [7:0]     TX_DATA_85_const_net_24;
wire   [7:0]     TX_DATA_86_const_net_24;
wire   [7:0]     TX_DATA_87_const_net_24;
wire   [7:0]     TX_DATA_88_const_net_24;
wire   [7:0]     TX_DATA_89_const_net_24;
wire   [7:0]     TX_DATA_90_const_net_24;
wire   [7:0]     TX_DATA_91_const_net_24;
wire   [7:0]     TX_DATA_92_const_net_24;
wire   [7:0]     TX_DATA_93_const_net_24;
wire   [7:0]     TX_DATA_94_const_net_24;
wire   [7:0]     TX_DATA_95_const_net_24;
wire   [7:0]     TX_DATA_96_const_net_24;
wire   [7:0]     TX_DATA_97_const_net_24;
wire   [7:0]     TX_DATA_98_const_net_24;
wire   [7:0]     TX_DATA_99_const_net_24;
wire   [7:0]     TX_DATA_100_const_net_24;
wire   [7:0]     TX_DATA_101_const_net_24;
wire   [7:0]     TX_DATA_102_const_net_24;
wire   [7:0]     TX_DATA_103_const_net_24;
wire   [7:0]     TX_DATA_104_const_net_24;
wire   [7:0]     TX_DATA_105_const_net_24;
wire   [7:0]     TX_DATA_106_const_net_24;
wire   [7:0]     TX_DATA_107_const_net_24;
wire   [7:0]     TX_DATA_108_const_net_24;
wire   [7:0]     TX_DATA_109_const_net_24;
wire   [7:0]     TX_DATA_110_const_net_24;
wire   [7:0]     TX_DATA_111_const_net_24;
wire   [7:0]     TX_DATA_112_const_net_24;
wire   [7:0]     TX_DATA_113_const_net_24;
wire   [7:0]     TX_DATA_114_const_net_24;
wire   [7:0]     TX_DATA_115_const_net_24;
wire   [7:0]     TX_DATA_116_const_net_24;
wire   [7:0]     TX_DATA_117_const_net_24;
wire   [7:0]     TX_DATA_118_const_net_24;
wire   [7:0]     TX_DATA_119_const_net_24;
wire   [7:0]     TX_DATA_120_const_net_24;
wire   [7:0]     TX_DATA_121_const_net_24;
wire   [7:0]     TX_DATA_122_const_net_24;
wire   [7:0]     TX_DATA_123_const_net_24;
wire   [7:0]     TX_DATA_124_const_net_24;
wire   [7:0]     TX_DATA_125_const_net_24;
wire   [7:0]     TX_DATA_126_const_net_24;
wire   [7:0]     TX_DATA_127_const_net_24;
wire   [3:0]     OE_DATA_1_const_net_22;
wire   [3:0]     OE_DATA_2_const_net_22;
wire   [3:0]     OE_DATA_3_const_net_22;
wire   [3:0]     OE_DATA_4_const_net_22;
wire   [3:0]     OE_DATA_5_const_net_22;
wire   [3:0]     OE_DATA_6_const_net_22;
wire   [3:0]     OE_DATA_7_const_net_22;
wire   [3:0]     OE_DATA_8_const_net_24;
wire   [3:0]     OE_DATA_9_const_net_24;
wire   [3:0]     OE_DATA_10_const_net_24;
wire   [3:0]     OE_DATA_11_const_net_24;
wire   [3:0]     OE_DATA_12_const_net_24;
wire   [3:0]     OE_DATA_13_const_net_24;
wire   [3:0]     OE_DATA_14_const_net_24;
wire   [3:0]     OE_DATA_15_const_net_24;
wire   [3:0]     OE_DATA_16_const_net_24;
wire   [3:0]     OE_DATA_17_const_net_24;
wire   [3:0]     OE_DATA_18_const_net_24;
wire   [3:0]     OE_DATA_19_const_net_24;
wire   [3:0]     OE_DATA_20_const_net_24;
wire   [3:0]     OE_DATA_21_const_net_24;
wire   [3:0]     OE_DATA_22_const_net_24;
wire   [3:0]     OE_DATA_23_const_net_24;
wire   [3:0]     OE_DATA_24_const_net_24;
wire   [3:0]     OE_DATA_25_const_net_24;
wire   [3:0]     OE_DATA_26_const_net_24;
wire   [3:0]     OE_DATA_27_const_net_24;
wire   [3:0]     OE_DATA_28_const_net_24;
wire   [3:0]     OE_DATA_29_const_net_24;
wire   [3:0]     OE_DATA_30_const_net_24;
wire   [3:0]     OE_DATA_31_const_net_24;
wire   [3:0]     OE_DATA_32_const_net_24;
wire   [3:0]     OE_DATA_33_const_net_24;
wire   [3:0]     OE_DATA_34_const_net_24;
wire   [3:0]     OE_DATA_35_const_net_24;
wire   [3:0]     OE_DATA_36_const_net_24;
wire   [3:0]     OE_DATA_37_const_net_24;
wire   [3:0]     OE_DATA_38_const_net_24;
wire   [3:0]     OE_DATA_39_const_net_24;
wire   [3:0]     OE_DATA_40_const_net_24;
wire   [3:0]     OE_DATA_41_const_net_24;
wire   [3:0]     OE_DATA_42_const_net_24;
wire   [3:0]     OE_DATA_43_const_net_24;
wire   [3:0]     OE_DATA_44_const_net_24;
wire   [3:0]     OE_DATA_45_const_net_24;
wire   [3:0]     OE_DATA_46_const_net_24;
wire   [3:0]     OE_DATA_47_const_net_24;
wire   [3:0]     OE_DATA_48_const_net_24;
wire   [3:0]     OE_DATA_49_const_net_24;
wire   [3:0]     OE_DATA_50_const_net_24;
wire   [3:0]     OE_DATA_51_const_net_24;
wire   [3:0]     OE_DATA_52_const_net_24;
wire   [3:0]     OE_DATA_53_const_net_24;
wire   [3:0]     OE_DATA_54_const_net_24;
wire   [3:0]     OE_DATA_55_const_net_24;
wire   [3:0]     OE_DATA_56_const_net_24;
wire   [3:0]     OE_DATA_57_const_net_24;
wire   [3:0]     OE_DATA_58_const_net_24;
wire   [3:0]     OE_DATA_59_const_net_24;
wire   [3:0]     OE_DATA_60_const_net_24;
wire   [3:0]     OE_DATA_61_const_net_24;
wire   [3:0]     OE_DATA_62_const_net_24;
wire   [3:0]     OE_DATA_63_const_net_24;
wire   [3:0]     OE_DATA_64_const_net_24;
wire   [3:0]     OE_DATA_65_const_net_24;
wire   [3:0]     OE_DATA_66_const_net_24;
wire   [3:0]     OE_DATA_67_const_net_24;
wire   [3:0]     OE_DATA_68_const_net_24;
wire   [3:0]     OE_DATA_69_const_net_24;
wire   [3:0]     OE_DATA_70_const_net_24;
wire   [3:0]     OE_DATA_71_const_net_24;
wire   [3:0]     OE_DATA_72_const_net_24;
wire   [3:0]     OE_DATA_73_const_net_24;
wire   [3:0]     OE_DATA_74_const_net_24;
wire   [3:0]     OE_DATA_75_const_net_24;
wire   [3:0]     OE_DATA_76_const_net_24;
wire   [3:0]     OE_DATA_77_const_net_24;
wire   [3:0]     OE_DATA_78_const_net_24;
wire   [3:0]     OE_DATA_79_const_net_24;
wire   [3:0]     OE_DATA_80_const_net_24;
wire   [3:0]     OE_DATA_81_const_net_24;
wire   [3:0]     OE_DATA_82_const_net_24;
wire   [3:0]     OE_DATA_83_const_net_24;
wire   [3:0]     OE_DATA_84_const_net_24;
wire   [3:0]     OE_DATA_85_const_net_24;
wire   [3:0]     OE_DATA_86_const_net_24;
wire   [3:0]     OE_DATA_87_const_net_24;
wire   [3:0]     OE_DATA_88_const_net_24;
wire   [3:0]     OE_DATA_89_const_net_24;
wire   [3:0]     OE_DATA_90_const_net_24;
wire   [3:0]     OE_DATA_91_const_net_24;
wire   [3:0]     OE_DATA_92_const_net_24;
wire   [3:0]     OE_DATA_93_const_net_24;
wire   [3:0]     OE_DATA_94_const_net_24;
wire   [3:0]     OE_DATA_95_const_net_24;
wire   [3:0]     OE_DATA_96_const_net_24;
wire   [3:0]     OE_DATA_97_const_net_24;
wire   [3:0]     OE_DATA_98_const_net_24;
wire   [3:0]     OE_DATA_99_const_net_24;
wire   [3:0]     OE_DATA_100_const_net_24;
wire   [3:0]     OE_DATA_101_const_net_24;
wire   [3:0]     OE_DATA_102_const_net_24;
wire   [3:0]     OE_DATA_103_const_net_24;
wire   [3:0]     OE_DATA_104_const_net_24;
wire   [3:0]     OE_DATA_105_const_net_24;
wire   [3:0]     OE_DATA_106_const_net_24;
wire   [3:0]     OE_DATA_107_const_net_24;
wire   [3:0]     OE_DATA_108_const_net_24;
wire   [3:0]     OE_DATA_109_const_net_24;
wire   [3:0]     OE_DATA_110_const_net_24;
wire   [3:0]     OE_DATA_111_const_net_24;
wire   [3:0]     OE_DATA_112_const_net_24;
wire   [3:0]     OE_DATA_113_const_net_24;
wire   [3:0]     OE_DATA_114_const_net_24;
wire   [3:0]     OE_DATA_115_const_net_24;
wire   [3:0]     OE_DATA_116_const_net_24;
wire   [3:0]     OE_DATA_117_const_net_24;
wire   [3:0]     OE_DATA_118_const_net_24;
wire   [3:0]     OE_DATA_119_const_net_24;
wire   [3:0]     OE_DATA_120_const_net_24;
wire   [3:0]     OE_DATA_121_const_net_24;
wire   [3:0]     OE_DATA_122_const_net_24;
wire   [3:0]     OE_DATA_123_const_net_24;
wire   [3:0]     OE_DATA_124_const_net_24;
wire   [3:0]     OE_DATA_125_const_net_24;
wire   [3:0]     OE_DATA_126_const_net_24;
wire   [3:0]     OE_DATA_127_const_net_24;
wire   [10:0]    CDR_CLK_B_SEL_const_net_2;
wire   [2:0]     FIFO_WR_PTR_const_net_19;
wire   [2:0]     FIFO_RD_PTR_const_net_19;
wire   [2:0]     EYE_MONITOR_LANE_WIDTH_const_net_21;
wire   [7:0]     TX_DATA_1_const_net_20;
wire   [7:0]     TX_DATA_2_const_net_22;
wire   [7:0]     TX_DATA_3_const_net_22;
wire   [7:0]     TX_DATA_4_const_net_22;
wire   [7:0]     TX_DATA_5_const_net_22;
wire   [7:0]     TX_DATA_6_const_net_22;
wire   [7:0]     TX_DATA_7_const_net_22;
wire   [7:0]     TX_DATA_8_const_net_24;
wire   [7:0]     TX_DATA_9_const_net_24;
wire   [7:0]     TX_DATA_10_const_net_24;
wire   [7:0]     TX_DATA_11_const_net_24;
wire   [7:0]     TX_DATA_12_const_net_25;
wire   [7:0]     TX_DATA_13_const_net_25;
wire   [7:0]     TX_DATA_14_const_net_25;
wire   [7:0]     TX_DATA_15_const_net_25;
wire   [7:0]     TX_DATA_16_const_net_25;
wire   [7:0]     TX_DATA_17_const_net_25;
wire   [7:0]     TX_DATA_18_const_net_25;
wire   [7:0]     TX_DATA_19_const_net_25;
wire   [7:0]     TX_DATA_20_const_net_25;
wire   [7:0]     TX_DATA_21_const_net_25;
wire   [7:0]     TX_DATA_22_const_net_25;
wire   [7:0]     TX_DATA_23_const_net_25;
wire   [7:0]     TX_DATA_24_const_net_25;
wire   [7:0]     TX_DATA_25_const_net_25;
wire   [7:0]     TX_DATA_26_const_net_25;
wire   [7:0]     TX_DATA_27_const_net_25;
wire   [7:0]     TX_DATA_28_const_net_25;
wire   [7:0]     TX_DATA_29_const_net_25;
wire   [7:0]     TX_DATA_30_const_net_25;
wire   [7:0]     TX_DATA_31_const_net_25;
wire   [7:0]     TX_DATA_32_const_net_25;
wire   [7:0]     TX_DATA_33_const_net_25;
wire   [7:0]     TX_DATA_34_const_net_25;
wire   [7:0]     TX_DATA_35_const_net_25;
wire   [7:0]     TX_DATA_36_const_net_25;
wire   [7:0]     TX_DATA_37_const_net_25;
wire   [7:0]     TX_DATA_38_const_net_25;
wire   [7:0]     TX_DATA_39_const_net_25;
wire   [7:0]     TX_DATA_40_const_net_25;
wire   [7:0]     TX_DATA_41_const_net_25;
wire   [7:0]     TX_DATA_42_const_net_25;
wire   [7:0]     TX_DATA_43_const_net_25;
wire   [7:0]     TX_DATA_44_const_net_25;
wire   [7:0]     TX_DATA_45_const_net_25;
wire   [7:0]     TX_DATA_46_const_net_25;
wire   [7:0]     TX_DATA_47_const_net_25;
wire   [7:0]     TX_DATA_48_const_net_25;
wire   [7:0]     TX_DATA_49_const_net_25;
wire   [7:0]     TX_DATA_50_const_net_25;
wire   [7:0]     TX_DATA_51_const_net_25;
wire   [7:0]     TX_DATA_52_const_net_25;
wire   [7:0]     TX_DATA_53_const_net_25;
wire   [7:0]     TX_DATA_54_const_net_25;
wire   [7:0]     TX_DATA_55_const_net_25;
wire   [7:0]     TX_DATA_56_const_net_25;
wire   [7:0]     TX_DATA_57_const_net_25;
wire   [7:0]     TX_DATA_58_const_net_25;
wire   [7:0]     TX_DATA_59_const_net_25;
wire   [7:0]     TX_DATA_60_const_net_25;
wire   [7:0]     TX_DATA_61_const_net_25;
wire   [7:0]     TX_DATA_62_const_net_25;
wire   [7:0]     TX_DATA_63_const_net_25;
wire   [7:0]     TX_DATA_64_const_net_25;
wire   [7:0]     TX_DATA_65_const_net_25;
wire   [7:0]     TX_DATA_66_const_net_25;
wire   [7:0]     TX_DATA_67_const_net_25;
wire   [7:0]     TX_DATA_68_const_net_25;
wire   [7:0]     TX_DATA_69_const_net_25;
wire   [7:0]     TX_DATA_70_const_net_25;
wire   [7:0]     TX_DATA_71_const_net_25;
wire   [7:0]     TX_DATA_72_const_net_25;
wire   [7:0]     TX_DATA_73_const_net_25;
wire   [7:0]     TX_DATA_74_const_net_25;
wire   [7:0]     TX_DATA_75_const_net_25;
wire   [7:0]     TX_DATA_76_const_net_25;
wire   [7:0]     TX_DATA_77_const_net_25;
wire   [7:0]     TX_DATA_78_const_net_25;
wire   [7:0]     TX_DATA_79_const_net_25;
wire   [7:0]     TX_DATA_80_const_net_25;
wire   [7:0]     TX_DATA_81_const_net_25;
wire   [7:0]     TX_DATA_82_const_net_25;
wire   [7:0]     TX_DATA_83_const_net_25;
wire   [7:0]     TX_DATA_84_const_net_25;
wire   [7:0]     TX_DATA_85_const_net_25;
wire   [7:0]     TX_DATA_86_const_net_25;
wire   [7:0]     TX_DATA_87_const_net_25;
wire   [7:0]     TX_DATA_88_const_net_25;
wire   [7:0]     TX_DATA_89_const_net_25;
wire   [7:0]     TX_DATA_90_const_net_25;
wire   [7:0]     TX_DATA_91_const_net_25;
wire   [7:0]     TX_DATA_92_const_net_25;
wire   [7:0]     TX_DATA_93_const_net_25;
wire   [7:0]     TX_DATA_94_const_net_25;
wire   [7:0]     TX_DATA_95_const_net_25;
wire   [7:0]     TX_DATA_96_const_net_25;
wire   [7:0]     TX_DATA_97_const_net_25;
wire   [7:0]     TX_DATA_98_const_net_25;
wire   [7:0]     TX_DATA_99_const_net_25;
wire   [7:0]     TX_DATA_100_const_net_25;
wire   [7:0]     TX_DATA_101_const_net_25;
wire   [7:0]     TX_DATA_102_const_net_25;
wire   [7:0]     TX_DATA_103_const_net_25;
wire   [7:0]     TX_DATA_104_const_net_25;
wire   [7:0]     TX_DATA_105_const_net_25;
wire   [7:0]     TX_DATA_106_const_net_25;
wire   [7:0]     TX_DATA_107_const_net_25;
wire   [7:0]     TX_DATA_108_const_net_25;
wire   [7:0]     TX_DATA_109_const_net_25;
wire   [7:0]     TX_DATA_110_const_net_25;
wire   [7:0]     TX_DATA_111_const_net_25;
wire   [7:0]     TX_DATA_112_const_net_25;
wire   [7:0]     TX_DATA_113_const_net_25;
wire   [7:0]     TX_DATA_114_const_net_25;
wire   [7:0]     TX_DATA_115_const_net_25;
wire   [7:0]     TX_DATA_116_const_net_25;
wire   [7:0]     TX_DATA_117_const_net_25;
wire   [7:0]     TX_DATA_118_const_net_25;
wire   [7:0]     TX_DATA_119_const_net_25;
wire   [7:0]     TX_DATA_120_const_net_25;
wire   [7:0]     TX_DATA_121_const_net_25;
wire   [7:0]     TX_DATA_122_const_net_25;
wire   [7:0]     TX_DATA_123_const_net_25;
wire   [7:0]     TX_DATA_124_const_net_25;
wire   [7:0]     TX_DATA_125_const_net_25;
wire   [7:0]     TX_DATA_126_const_net_25;
wire   [7:0]     TX_DATA_127_const_net_25;
wire   [3:0]     OE_DATA_1_const_net_23;
wire   [3:0]     OE_DATA_2_const_net_23;
wire   [3:0]     OE_DATA_3_const_net_23;
wire   [3:0]     OE_DATA_4_const_net_23;
wire   [3:0]     OE_DATA_5_const_net_23;
wire   [3:0]     OE_DATA_6_const_net_23;
wire   [3:0]     OE_DATA_7_const_net_23;
wire   [3:0]     OE_DATA_8_const_net_25;
wire   [3:0]     OE_DATA_9_const_net_25;
wire   [3:0]     OE_DATA_10_const_net_25;
wire   [3:0]     OE_DATA_11_const_net_25;
wire   [3:0]     OE_DATA_12_const_net_25;
wire   [3:0]     OE_DATA_13_const_net_25;
wire   [3:0]     OE_DATA_14_const_net_25;
wire   [3:0]     OE_DATA_15_const_net_25;
wire   [3:0]     OE_DATA_16_const_net_25;
wire   [3:0]     OE_DATA_17_const_net_25;
wire   [3:0]     OE_DATA_18_const_net_25;
wire   [3:0]     OE_DATA_19_const_net_25;
wire   [3:0]     OE_DATA_20_const_net_25;
wire   [3:0]     OE_DATA_21_const_net_25;
wire   [3:0]     OE_DATA_22_const_net_25;
wire   [3:0]     OE_DATA_23_const_net_25;
wire   [3:0]     OE_DATA_24_const_net_25;
wire   [3:0]     OE_DATA_25_const_net_25;
wire   [3:0]     OE_DATA_26_const_net_25;
wire   [3:0]     OE_DATA_27_const_net_25;
wire   [3:0]     OE_DATA_28_const_net_25;
wire   [3:0]     OE_DATA_29_const_net_25;
wire   [3:0]     OE_DATA_30_const_net_25;
wire   [3:0]     OE_DATA_31_const_net_25;
wire   [3:0]     OE_DATA_32_const_net_25;
wire   [3:0]     OE_DATA_33_const_net_25;
wire   [3:0]     OE_DATA_34_const_net_25;
wire   [3:0]     OE_DATA_35_const_net_25;
wire   [3:0]     OE_DATA_36_const_net_25;
wire   [3:0]     OE_DATA_37_const_net_25;
wire   [3:0]     OE_DATA_38_const_net_25;
wire   [3:0]     OE_DATA_39_const_net_25;
wire   [3:0]     OE_DATA_40_const_net_25;
wire   [3:0]     OE_DATA_41_const_net_25;
wire   [3:0]     OE_DATA_42_const_net_25;
wire   [3:0]     OE_DATA_43_const_net_25;
wire   [3:0]     OE_DATA_44_const_net_25;
wire   [3:0]     OE_DATA_45_const_net_25;
wire   [3:0]     OE_DATA_46_const_net_25;
wire   [3:0]     OE_DATA_47_const_net_25;
wire   [3:0]     OE_DATA_48_const_net_25;
wire   [3:0]     OE_DATA_49_const_net_25;
wire   [3:0]     OE_DATA_50_const_net_25;
wire   [3:0]     OE_DATA_51_const_net_25;
wire   [3:0]     OE_DATA_52_const_net_25;
wire   [3:0]     OE_DATA_53_const_net_25;
wire   [3:0]     OE_DATA_54_const_net_25;
wire   [3:0]     OE_DATA_55_const_net_25;
wire   [3:0]     OE_DATA_56_const_net_25;
wire   [3:0]     OE_DATA_57_const_net_25;
wire   [3:0]     OE_DATA_58_const_net_25;
wire   [3:0]     OE_DATA_59_const_net_25;
wire   [3:0]     OE_DATA_60_const_net_25;
wire   [3:0]     OE_DATA_61_const_net_25;
wire   [3:0]     OE_DATA_62_const_net_25;
wire   [3:0]     OE_DATA_63_const_net_25;
wire   [3:0]     OE_DATA_64_const_net_25;
wire   [3:0]     OE_DATA_65_const_net_25;
wire   [3:0]     OE_DATA_66_const_net_25;
wire   [3:0]     OE_DATA_67_const_net_25;
wire   [3:0]     OE_DATA_68_const_net_25;
wire   [3:0]     OE_DATA_69_const_net_25;
wire   [3:0]     OE_DATA_70_const_net_25;
wire   [3:0]     OE_DATA_71_const_net_25;
wire   [3:0]     OE_DATA_72_const_net_25;
wire   [3:0]     OE_DATA_73_const_net_25;
wire   [3:0]     OE_DATA_74_const_net_25;
wire   [3:0]     OE_DATA_75_const_net_25;
wire   [3:0]     OE_DATA_76_const_net_25;
wire   [3:0]     OE_DATA_77_const_net_25;
wire   [3:0]     OE_DATA_78_const_net_25;
wire   [3:0]     OE_DATA_79_const_net_25;
wire   [3:0]     OE_DATA_80_const_net_25;
wire   [3:0]     OE_DATA_81_const_net_25;
wire   [3:0]     OE_DATA_82_const_net_25;
wire   [3:0]     OE_DATA_83_const_net_25;
wire   [3:0]     OE_DATA_84_const_net_25;
wire   [3:0]     OE_DATA_85_const_net_25;
wire   [3:0]     OE_DATA_86_const_net_25;
wire   [3:0]     OE_DATA_87_const_net_25;
wire   [3:0]     OE_DATA_88_const_net_25;
wire   [3:0]     OE_DATA_89_const_net_25;
wire   [3:0]     OE_DATA_90_const_net_25;
wire   [3:0]     OE_DATA_91_const_net_25;
wire   [3:0]     OE_DATA_92_const_net_25;
wire   [3:0]     OE_DATA_93_const_net_25;
wire   [3:0]     OE_DATA_94_const_net_25;
wire   [3:0]     OE_DATA_95_const_net_25;
wire   [3:0]     OE_DATA_96_const_net_25;
wire   [3:0]     OE_DATA_97_const_net_25;
wire   [3:0]     OE_DATA_98_const_net_25;
wire   [3:0]     OE_DATA_99_const_net_25;
wire   [3:0]     OE_DATA_100_const_net_25;
wire   [3:0]     OE_DATA_101_const_net_25;
wire   [3:0]     OE_DATA_102_const_net_25;
wire   [3:0]     OE_DATA_103_const_net_25;
wire   [3:0]     OE_DATA_104_const_net_25;
wire   [3:0]     OE_DATA_105_const_net_25;
wire   [3:0]     OE_DATA_106_const_net_25;
wire   [3:0]     OE_DATA_107_const_net_25;
wire   [3:0]     OE_DATA_108_const_net_25;
wire   [3:0]     OE_DATA_109_const_net_25;
wire   [3:0]     OE_DATA_110_const_net_25;
wire   [3:0]     OE_DATA_111_const_net_25;
wire   [3:0]     OE_DATA_112_const_net_25;
wire   [3:0]     OE_DATA_113_const_net_25;
wire   [3:0]     OE_DATA_114_const_net_25;
wire   [3:0]     OE_DATA_115_const_net_25;
wire   [3:0]     OE_DATA_116_const_net_25;
wire   [3:0]     OE_DATA_117_const_net_25;
wire   [3:0]     OE_DATA_118_const_net_25;
wire   [3:0]     OE_DATA_119_const_net_25;
wire   [3:0]     OE_DATA_120_const_net_25;
wire   [3:0]     OE_DATA_121_const_net_25;
wire   [3:0]     OE_DATA_122_const_net_25;
wire   [3:0]     OE_DATA_123_const_net_25;
wire   [3:0]     OE_DATA_124_const_net_25;
wire   [3:0]     OE_DATA_125_const_net_25;
wire   [3:0]     OE_DATA_126_const_net_25;
wire   [3:0]     OE_DATA_127_const_net_25;
wire   [7:0]     TX_DATA_8_const_net_25;
wire   [7:0]     TX_DATA_9_const_net_25;
wire   [7:0]     TX_DATA_10_const_net_25;
wire   [7:0]     TX_DATA_11_const_net_25;
wire   [7:0]     TX_DATA_12_const_net_26;
wire   [7:0]     TX_DATA_13_const_net_26;
wire   [7:0]     TX_DATA_14_const_net_26;
wire   [7:0]     TX_DATA_15_const_net_26;
wire   [7:0]     TX_DATA_16_const_net_26;
wire   [7:0]     TX_DATA_17_const_net_26;
wire   [7:0]     TX_DATA_18_const_net_26;
wire   [7:0]     TX_DATA_19_const_net_26;
wire   [7:0]     TX_DATA_20_const_net_26;
wire   [7:0]     TX_DATA_21_const_net_26;
wire   [7:0]     TX_DATA_22_const_net_26;
wire   [7:0]     TX_DATA_23_const_net_26;
wire   [7:0]     TX_DATA_24_const_net_26;
wire   [7:0]     TX_DATA_25_const_net_26;
wire   [7:0]     TX_DATA_26_const_net_26;
wire   [7:0]     TX_DATA_27_const_net_26;
wire   [7:0]     TX_DATA_28_const_net_26;
wire   [7:0]     TX_DATA_29_const_net_26;
wire   [7:0]     TX_DATA_30_const_net_26;
wire   [7:0]     TX_DATA_31_const_net_26;
wire   [7:0]     TX_DATA_32_const_net_26;
wire   [7:0]     TX_DATA_33_const_net_26;
wire   [7:0]     TX_DATA_34_const_net_26;
wire   [7:0]     TX_DATA_35_const_net_26;
wire   [7:0]     TX_DATA_36_const_net_26;
wire   [7:0]     TX_DATA_37_const_net_26;
wire   [7:0]     TX_DATA_38_const_net_26;
wire   [7:0]     TX_DATA_39_const_net_26;
wire   [7:0]     TX_DATA_40_const_net_26;
wire   [7:0]     TX_DATA_41_const_net_26;
wire   [7:0]     TX_DATA_42_const_net_26;
wire   [7:0]     TX_DATA_43_const_net_26;
wire   [7:0]     TX_DATA_44_const_net_26;
wire   [7:0]     TX_DATA_45_const_net_26;
wire   [7:0]     TX_DATA_46_const_net_26;
wire   [7:0]     TX_DATA_47_const_net_26;
wire   [7:0]     TX_DATA_48_const_net_26;
wire   [7:0]     TX_DATA_49_const_net_26;
wire   [7:0]     TX_DATA_50_const_net_26;
wire   [7:0]     TX_DATA_51_const_net_26;
wire   [7:0]     TX_DATA_52_const_net_26;
wire   [7:0]     TX_DATA_53_const_net_26;
wire   [7:0]     TX_DATA_54_const_net_26;
wire   [7:0]     TX_DATA_55_const_net_26;
wire   [7:0]     TX_DATA_56_const_net_26;
wire   [7:0]     TX_DATA_57_const_net_26;
wire   [7:0]     TX_DATA_58_const_net_26;
wire   [7:0]     TX_DATA_59_const_net_26;
wire   [7:0]     TX_DATA_60_const_net_26;
wire   [7:0]     TX_DATA_61_const_net_26;
wire   [7:0]     TX_DATA_62_const_net_26;
wire   [7:0]     TX_DATA_63_const_net_26;
wire   [7:0]     TX_DATA_64_const_net_26;
wire   [7:0]     TX_DATA_65_const_net_26;
wire   [7:0]     TX_DATA_66_const_net_26;
wire   [7:0]     TX_DATA_67_const_net_26;
wire   [7:0]     TX_DATA_68_const_net_26;
wire   [7:0]     TX_DATA_69_const_net_26;
wire   [7:0]     TX_DATA_70_const_net_26;
wire   [7:0]     TX_DATA_71_const_net_26;
wire   [7:0]     TX_DATA_72_const_net_26;
wire   [7:0]     TX_DATA_73_const_net_26;
wire   [7:0]     TX_DATA_74_const_net_26;
wire   [7:0]     TX_DATA_75_const_net_26;
wire   [7:0]     TX_DATA_76_const_net_26;
wire   [7:0]     TX_DATA_77_const_net_26;
wire   [7:0]     TX_DATA_78_const_net_26;
wire   [7:0]     TX_DATA_79_const_net_26;
wire   [7:0]     TX_DATA_80_const_net_26;
wire   [7:0]     TX_DATA_81_const_net_26;
wire   [7:0]     TX_DATA_82_const_net_26;
wire   [7:0]     TX_DATA_83_const_net_26;
wire   [7:0]     TX_DATA_84_const_net_26;
wire   [7:0]     TX_DATA_85_const_net_26;
wire   [7:0]     TX_DATA_86_const_net_26;
wire   [7:0]     TX_DATA_87_const_net_26;
wire   [7:0]     TX_DATA_88_const_net_26;
wire   [7:0]     TX_DATA_89_const_net_26;
wire   [7:0]     TX_DATA_90_const_net_26;
wire   [7:0]     TX_DATA_91_const_net_26;
wire   [7:0]     TX_DATA_92_const_net_26;
wire   [7:0]     TX_DATA_93_const_net_26;
wire   [7:0]     TX_DATA_94_const_net_26;
wire   [7:0]     TX_DATA_95_const_net_26;
wire   [7:0]     TX_DATA_96_const_net_26;
wire   [7:0]     TX_DATA_97_const_net_26;
wire   [7:0]     TX_DATA_98_const_net_26;
wire   [7:0]     TX_DATA_99_const_net_26;
wire   [7:0]     TX_DATA_100_const_net_26;
wire   [7:0]     TX_DATA_101_const_net_26;
wire   [7:0]     TX_DATA_102_const_net_26;
wire   [7:0]     TX_DATA_103_const_net_26;
wire   [7:0]     TX_DATA_104_const_net_26;
wire   [7:0]     TX_DATA_105_const_net_26;
wire   [7:0]     TX_DATA_106_const_net_26;
wire   [7:0]     TX_DATA_107_const_net_26;
wire   [7:0]     TX_DATA_108_const_net_26;
wire   [7:0]     TX_DATA_109_const_net_26;
wire   [7:0]     TX_DATA_110_const_net_26;
wire   [7:0]     TX_DATA_111_const_net_26;
wire   [7:0]     TX_DATA_112_const_net_26;
wire   [7:0]     TX_DATA_113_const_net_26;
wire   [7:0]     TX_DATA_114_const_net_26;
wire   [7:0]     TX_DATA_115_const_net_26;
wire   [7:0]     TX_DATA_116_const_net_26;
wire   [7:0]     TX_DATA_117_const_net_26;
wire   [7:0]     TX_DATA_118_const_net_26;
wire   [7:0]     TX_DATA_119_const_net_26;
wire   [7:0]     TX_DATA_120_const_net_26;
wire   [7:0]     TX_DATA_121_const_net_26;
wire   [7:0]     TX_DATA_122_const_net_26;
wire   [7:0]     TX_DATA_123_const_net_26;
wire   [7:0]     TX_DATA_124_const_net_26;
wire   [7:0]     TX_DATA_125_const_net_26;
wire   [7:0]     TX_DATA_126_const_net_26;
wire   [7:0]     TX_DATA_127_const_net_26;
wire   [3:0]     OE_DATA_8_const_net_26;
wire   [3:0]     OE_DATA_9_const_net_26;
wire   [3:0]     OE_DATA_10_const_net_26;
wire   [3:0]     OE_DATA_11_const_net_26;
wire   [3:0]     OE_DATA_12_const_net_26;
wire   [3:0]     OE_DATA_13_const_net_26;
wire   [3:0]     OE_DATA_14_const_net_26;
wire   [3:0]     OE_DATA_15_const_net_26;
wire   [3:0]     OE_DATA_16_const_net_26;
wire   [3:0]     OE_DATA_17_const_net_26;
wire   [3:0]     OE_DATA_18_const_net_26;
wire   [3:0]     OE_DATA_19_const_net_26;
wire   [3:0]     OE_DATA_20_const_net_26;
wire   [3:0]     OE_DATA_21_const_net_26;
wire   [3:0]     OE_DATA_22_const_net_26;
wire   [3:0]     OE_DATA_23_const_net_26;
wire   [3:0]     OE_DATA_24_const_net_26;
wire   [3:0]     OE_DATA_25_const_net_26;
wire   [3:0]     OE_DATA_26_const_net_26;
wire   [3:0]     OE_DATA_27_const_net_26;
wire   [3:0]     OE_DATA_28_const_net_26;
wire   [3:0]     OE_DATA_29_const_net_26;
wire   [3:0]     OE_DATA_30_const_net_26;
wire   [3:0]     OE_DATA_31_const_net_26;
wire   [3:0]     OE_DATA_32_const_net_26;
wire   [3:0]     OE_DATA_33_const_net_26;
wire   [3:0]     OE_DATA_34_const_net_26;
wire   [3:0]     OE_DATA_35_const_net_26;
wire   [3:0]     OE_DATA_36_const_net_26;
wire   [3:0]     OE_DATA_37_const_net_26;
wire   [3:0]     OE_DATA_38_const_net_26;
wire   [3:0]     OE_DATA_39_const_net_26;
wire   [3:0]     OE_DATA_40_const_net_26;
wire   [3:0]     OE_DATA_41_const_net_26;
wire   [3:0]     OE_DATA_42_const_net_26;
wire   [3:0]     OE_DATA_43_const_net_26;
wire   [3:0]     OE_DATA_44_const_net_26;
wire   [3:0]     OE_DATA_45_const_net_26;
wire   [3:0]     OE_DATA_46_const_net_26;
wire   [3:0]     OE_DATA_47_const_net_26;
wire   [3:0]     OE_DATA_48_const_net_26;
wire   [3:0]     OE_DATA_49_const_net_26;
wire   [3:0]     OE_DATA_50_const_net_26;
wire   [3:0]     OE_DATA_51_const_net_26;
wire   [3:0]     OE_DATA_52_const_net_26;
wire   [3:0]     OE_DATA_53_const_net_26;
wire   [3:0]     OE_DATA_54_const_net_26;
wire   [3:0]     OE_DATA_55_const_net_26;
wire   [3:0]     OE_DATA_56_const_net_26;
wire   [3:0]     OE_DATA_57_const_net_26;
wire   [3:0]     OE_DATA_58_const_net_26;
wire   [3:0]     OE_DATA_59_const_net_26;
wire   [3:0]     OE_DATA_60_const_net_26;
wire   [3:0]     OE_DATA_61_const_net_26;
wire   [3:0]     OE_DATA_62_const_net_26;
wire   [3:0]     OE_DATA_63_const_net_26;
wire   [3:0]     OE_DATA_64_const_net_26;
wire   [3:0]     OE_DATA_65_const_net_26;
wire   [3:0]     OE_DATA_66_const_net_26;
wire   [3:0]     OE_DATA_67_const_net_26;
wire   [3:0]     OE_DATA_68_const_net_26;
wire   [3:0]     OE_DATA_69_const_net_26;
wire   [3:0]     OE_DATA_70_const_net_26;
wire   [3:0]     OE_DATA_71_const_net_26;
wire   [3:0]     OE_DATA_72_const_net_26;
wire   [3:0]     OE_DATA_73_const_net_26;
wire   [3:0]     OE_DATA_74_const_net_26;
wire   [3:0]     OE_DATA_75_const_net_26;
wire   [3:0]     OE_DATA_76_const_net_26;
wire   [3:0]     OE_DATA_77_const_net_26;
wire   [3:0]     OE_DATA_78_const_net_26;
wire   [3:0]     OE_DATA_79_const_net_26;
wire   [3:0]     OE_DATA_80_const_net_26;
wire   [3:0]     OE_DATA_81_const_net_26;
wire   [3:0]     OE_DATA_82_const_net_26;
wire   [3:0]     OE_DATA_83_const_net_26;
wire   [3:0]     OE_DATA_84_const_net_26;
wire   [3:0]     OE_DATA_85_const_net_26;
wire   [3:0]     OE_DATA_86_const_net_26;
wire   [3:0]     OE_DATA_87_const_net_26;
wire   [3:0]     OE_DATA_88_const_net_26;
wire   [3:0]     OE_DATA_89_const_net_26;
wire   [3:0]     OE_DATA_90_const_net_26;
wire   [3:0]     OE_DATA_91_const_net_26;
wire   [3:0]     OE_DATA_92_const_net_26;
wire   [3:0]     OE_DATA_93_const_net_26;
wire   [3:0]     OE_DATA_94_const_net_26;
wire   [3:0]     OE_DATA_95_const_net_26;
wire   [3:0]     OE_DATA_96_const_net_26;
wire   [3:0]     OE_DATA_97_const_net_26;
wire   [3:0]     OE_DATA_98_const_net_26;
wire   [3:0]     OE_DATA_99_const_net_26;
wire   [3:0]     OE_DATA_100_const_net_26;
wire   [3:0]     OE_DATA_101_const_net_26;
wire   [3:0]     OE_DATA_102_const_net_26;
wire   [3:0]     OE_DATA_103_const_net_26;
wire   [3:0]     OE_DATA_104_const_net_26;
wire   [3:0]     OE_DATA_105_const_net_26;
wire   [3:0]     OE_DATA_106_const_net_26;
wire   [3:0]     OE_DATA_107_const_net_26;
wire   [3:0]     OE_DATA_108_const_net_26;
wire   [3:0]     OE_DATA_109_const_net_26;
wire   [3:0]     OE_DATA_110_const_net_26;
wire   [3:0]     OE_DATA_111_const_net_26;
wire   [3:0]     OE_DATA_112_const_net_26;
wire   [3:0]     OE_DATA_113_const_net_26;
wire   [3:0]     OE_DATA_114_const_net_26;
wire   [3:0]     OE_DATA_115_const_net_26;
wire   [3:0]     OE_DATA_116_const_net_26;
wire   [3:0]     OE_DATA_117_const_net_26;
wire   [3:0]     OE_DATA_118_const_net_26;
wire   [3:0]     OE_DATA_119_const_net_26;
wire   [3:0]     OE_DATA_120_const_net_26;
wire   [3:0]     OE_DATA_121_const_net_26;
wire   [3:0]     OE_DATA_122_const_net_26;
wire   [3:0]     OE_DATA_123_const_net_26;
wire   [3:0]     OE_DATA_124_const_net_26;
wire   [3:0]     OE_DATA_125_const_net_26;
wire   [3:0]     OE_DATA_126_const_net_26;
wire   [3:0]     OE_DATA_127_const_net_26;
wire   [7:0]     PAD_I_const_net_5;
wire   [7:0]     PAD_N_const_net_5;
wire   [7:0]     PAD_I_N_const_net_5;
wire   [7:0]     TX_DATA_1_const_net_21;
wire   [7:0]     TX_DATA_2_const_net_23;
wire   [7:0]     TX_DATA_3_const_net_23;
wire   [7:0]     TX_DATA_4_const_net_23;
wire   [7:0]     TX_DATA_5_const_net_23;
wire   [7:0]     TX_DATA_6_const_net_23;
wire   [7:0]     TX_DATA_7_const_net_23;
wire   [7:0]     TX_DATA_8_const_net_26;
wire   [7:0]     TX_DATA_9_const_net_26;
wire   [7:0]     TX_DATA_10_const_net_26;
wire   [7:0]     TX_DATA_11_const_net_26;
wire   [7:0]     TX_DATA_12_const_net_27;
wire   [7:0]     TX_DATA_13_const_net_27;
wire   [7:0]     TX_DATA_14_const_net_27;
wire   [7:0]     TX_DATA_15_const_net_27;
wire   [7:0]     TX_DATA_16_const_net_27;
wire   [7:0]     TX_DATA_17_const_net_27;
wire   [7:0]     TX_DATA_18_const_net_27;
wire   [7:0]     TX_DATA_19_const_net_27;
wire   [7:0]     TX_DATA_20_const_net_27;
wire   [7:0]     TX_DATA_21_const_net_27;
wire   [7:0]     TX_DATA_22_const_net_27;
wire   [7:0]     TX_DATA_23_const_net_27;
wire   [7:0]     TX_DATA_24_const_net_27;
wire   [7:0]     TX_DATA_25_const_net_27;
wire   [7:0]     TX_DATA_26_const_net_27;
wire   [7:0]     TX_DATA_27_const_net_27;
wire   [7:0]     TX_DATA_28_const_net_27;
wire   [7:0]     TX_DATA_29_const_net_27;
wire   [7:0]     TX_DATA_30_const_net_27;
wire   [7:0]     TX_DATA_31_const_net_27;
wire   [7:0]     TX_DATA_32_const_net_27;
wire   [7:0]     TX_DATA_33_const_net_27;
wire   [7:0]     TX_DATA_34_const_net_27;
wire   [7:0]     TX_DATA_35_const_net_27;
wire   [7:0]     TX_DATA_36_const_net_27;
wire   [7:0]     TX_DATA_37_const_net_27;
wire   [7:0]     TX_DATA_38_const_net_27;
wire   [7:0]     TX_DATA_39_const_net_27;
wire   [7:0]     TX_DATA_40_const_net_27;
wire   [7:0]     TX_DATA_41_const_net_27;
wire   [7:0]     TX_DATA_42_const_net_27;
wire   [7:0]     TX_DATA_43_const_net_27;
wire   [7:0]     TX_DATA_44_const_net_27;
wire   [7:0]     TX_DATA_45_const_net_27;
wire   [7:0]     TX_DATA_46_const_net_27;
wire   [7:0]     TX_DATA_47_const_net_27;
wire   [7:0]     TX_DATA_48_const_net_27;
wire   [7:0]     TX_DATA_49_const_net_27;
wire   [7:0]     TX_DATA_50_const_net_27;
wire   [7:0]     TX_DATA_51_const_net_27;
wire   [7:0]     TX_DATA_52_const_net_27;
wire   [7:0]     TX_DATA_53_const_net_27;
wire   [7:0]     TX_DATA_54_const_net_27;
wire   [7:0]     TX_DATA_55_const_net_27;
wire   [7:0]     TX_DATA_56_const_net_27;
wire   [7:0]     TX_DATA_57_const_net_27;
wire   [7:0]     TX_DATA_58_const_net_27;
wire   [7:0]     TX_DATA_59_const_net_27;
wire   [7:0]     TX_DATA_60_const_net_27;
wire   [7:0]     TX_DATA_61_const_net_27;
wire   [7:0]     TX_DATA_62_const_net_27;
wire   [7:0]     TX_DATA_63_const_net_27;
wire   [7:0]     TX_DATA_64_const_net_27;
wire   [7:0]     TX_DATA_65_const_net_27;
wire   [7:0]     TX_DATA_66_const_net_27;
wire   [7:0]     TX_DATA_67_const_net_27;
wire   [7:0]     TX_DATA_68_const_net_27;
wire   [7:0]     TX_DATA_69_const_net_27;
wire   [7:0]     TX_DATA_70_const_net_27;
wire   [7:0]     TX_DATA_71_const_net_27;
wire   [7:0]     TX_DATA_72_const_net_27;
wire   [7:0]     TX_DATA_73_const_net_27;
wire   [7:0]     TX_DATA_74_const_net_27;
wire   [7:0]     TX_DATA_75_const_net_27;
wire   [7:0]     TX_DATA_76_const_net_27;
wire   [7:0]     TX_DATA_77_const_net_27;
wire   [7:0]     TX_DATA_78_const_net_27;
wire   [7:0]     TX_DATA_79_const_net_27;
wire   [7:0]     TX_DATA_80_const_net_27;
wire   [7:0]     TX_DATA_81_const_net_27;
wire   [7:0]     TX_DATA_82_const_net_27;
wire   [7:0]     TX_DATA_83_const_net_27;
wire   [7:0]     TX_DATA_84_const_net_27;
wire   [7:0]     TX_DATA_85_const_net_27;
wire   [7:0]     TX_DATA_86_const_net_27;
wire   [7:0]     TX_DATA_87_const_net_27;
wire   [7:0]     TX_DATA_88_const_net_27;
wire   [7:0]     TX_DATA_89_const_net_27;
wire   [7:0]     TX_DATA_90_const_net_27;
wire   [7:0]     TX_DATA_91_const_net_27;
wire   [7:0]     TX_DATA_92_const_net_27;
wire   [7:0]     TX_DATA_93_const_net_27;
wire   [7:0]     TX_DATA_94_const_net_27;
wire   [7:0]     TX_DATA_95_const_net_27;
wire   [7:0]     TX_DATA_96_const_net_27;
wire   [7:0]     TX_DATA_97_const_net_27;
wire   [7:0]     TX_DATA_98_const_net_27;
wire   [7:0]     TX_DATA_99_const_net_27;
wire   [7:0]     TX_DATA_100_const_net_27;
wire   [7:0]     TX_DATA_101_const_net_27;
wire   [7:0]     TX_DATA_102_const_net_27;
wire   [7:0]     TX_DATA_103_const_net_27;
wire   [7:0]     TX_DATA_104_const_net_27;
wire   [7:0]     TX_DATA_105_const_net_27;
wire   [7:0]     TX_DATA_106_const_net_27;
wire   [7:0]     TX_DATA_107_const_net_27;
wire   [7:0]     TX_DATA_108_const_net_27;
wire   [7:0]     TX_DATA_109_const_net_27;
wire   [7:0]     TX_DATA_110_const_net_27;
wire   [7:0]     TX_DATA_111_const_net_27;
wire   [7:0]     TX_DATA_112_const_net_27;
wire   [7:0]     TX_DATA_113_const_net_27;
wire   [7:0]     TX_DATA_114_const_net_27;
wire   [7:0]     TX_DATA_115_const_net_27;
wire   [7:0]     TX_DATA_116_const_net_27;
wire   [7:0]     TX_DATA_117_const_net_27;
wire   [7:0]     TX_DATA_118_const_net_27;
wire   [7:0]     TX_DATA_119_const_net_27;
wire   [7:0]     TX_DATA_120_const_net_27;
wire   [7:0]     TX_DATA_121_const_net_27;
wire   [7:0]     TX_DATA_122_const_net_27;
wire   [7:0]     TX_DATA_123_const_net_27;
wire   [7:0]     TX_DATA_124_const_net_27;
wire   [7:0]     TX_DATA_125_const_net_27;
wire   [7:0]     TX_DATA_126_const_net_27;
wire   [7:0]     TX_DATA_127_const_net_27;
wire   [3:0]     OE_DATA_1_const_net_24;
wire   [3:0]     OE_DATA_2_const_net_24;
wire   [3:0]     OE_DATA_3_const_net_24;
wire   [3:0]     OE_DATA_4_const_net_24;
wire   [3:0]     OE_DATA_5_const_net_24;
wire   [3:0]     OE_DATA_6_const_net_24;
wire   [3:0]     OE_DATA_7_const_net_24;
wire   [3:0]     OE_DATA_8_const_net_27;
wire   [3:0]     OE_DATA_9_const_net_27;
wire   [3:0]     OE_DATA_10_const_net_27;
wire   [3:0]     OE_DATA_11_const_net_27;
wire   [3:0]     OE_DATA_12_const_net_27;
wire   [3:0]     OE_DATA_13_const_net_27;
wire   [3:0]     OE_DATA_14_const_net_27;
wire   [3:0]     OE_DATA_15_const_net_27;
wire   [3:0]     OE_DATA_16_const_net_27;
wire   [3:0]     OE_DATA_17_const_net_27;
wire   [3:0]     OE_DATA_18_const_net_27;
wire   [3:0]     OE_DATA_19_const_net_27;
wire   [3:0]     OE_DATA_20_const_net_27;
wire   [3:0]     OE_DATA_21_const_net_27;
wire   [3:0]     OE_DATA_22_const_net_27;
wire   [3:0]     OE_DATA_23_const_net_27;
wire   [3:0]     OE_DATA_24_const_net_27;
wire   [3:0]     OE_DATA_25_const_net_27;
wire   [3:0]     OE_DATA_26_const_net_27;
wire   [3:0]     OE_DATA_27_const_net_27;
wire   [3:0]     OE_DATA_28_const_net_27;
wire   [3:0]     OE_DATA_29_const_net_27;
wire   [3:0]     OE_DATA_30_const_net_27;
wire   [3:0]     OE_DATA_31_const_net_27;
wire   [3:0]     OE_DATA_32_const_net_27;
wire   [3:0]     OE_DATA_33_const_net_27;
wire   [3:0]     OE_DATA_34_const_net_27;
wire   [3:0]     OE_DATA_35_const_net_27;
wire   [3:0]     OE_DATA_36_const_net_27;
wire   [3:0]     OE_DATA_37_const_net_27;
wire   [3:0]     OE_DATA_38_const_net_27;
wire   [3:0]     OE_DATA_39_const_net_27;
wire   [3:0]     OE_DATA_40_const_net_27;
wire   [3:0]     OE_DATA_41_const_net_27;
wire   [3:0]     OE_DATA_42_const_net_27;
wire   [3:0]     OE_DATA_43_const_net_27;
wire   [3:0]     OE_DATA_44_const_net_27;
wire   [3:0]     OE_DATA_45_const_net_27;
wire   [3:0]     OE_DATA_46_const_net_27;
wire   [3:0]     OE_DATA_47_const_net_27;
wire   [3:0]     OE_DATA_48_const_net_27;
wire   [3:0]     OE_DATA_49_const_net_27;
wire   [3:0]     OE_DATA_50_const_net_27;
wire   [3:0]     OE_DATA_51_const_net_27;
wire   [3:0]     OE_DATA_52_const_net_27;
wire   [3:0]     OE_DATA_53_const_net_27;
wire   [3:0]     OE_DATA_54_const_net_27;
wire   [3:0]     OE_DATA_55_const_net_27;
wire   [3:0]     OE_DATA_56_const_net_27;
wire   [3:0]     OE_DATA_57_const_net_27;
wire   [3:0]     OE_DATA_58_const_net_27;
wire   [3:0]     OE_DATA_59_const_net_27;
wire   [3:0]     OE_DATA_60_const_net_27;
wire   [3:0]     OE_DATA_61_const_net_27;
wire   [3:0]     OE_DATA_62_const_net_27;
wire   [3:0]     OE_DATA_63_const_net_27;
wire   [3:0]     OE_DATA_64_const_net_27;
wire   [3:0]     OE_DATA_65_const_net_27;
wire   [3:0]     OE_DATA_66_const_net_27;
wire   [3:0]     OE_DATA_67_const_net_27;
wire   [3:0]     OE_DATA_68_const_net_27;
wire   [3:0]     OE_DATA_69_const_net_27;
wire   [3:0]     OE_DATA_70_const_net_27;
wire   [3:0]     OE_DATA_71_const_net_27;
wire   [3:0]     OE_DATA_72_const_net_27;
wire   [3:0]     OE_DATA_73_const_net_27;
wire   [3:0]     OE_DATA_74_const_net_27;
wire   [3:0]     OE_DATA_75_const_net_27;
wire   [3:0]     OE_DATA_76_const_net_27;
wire   [3:0]     OE_DATA_77_const_net_27;
wire   [3:0]     OE_DATA_78_const_net_27;
wire   [3:0]     OE_DATA_79_const_net_27;
wire   [3:0]     OE_DATA_80_const_net_27;
wire   [3:0]     OE_DATA_81_const_net_27;
wire   [3:0]     OE_DATA_82_const_net_27;
wire   [3:0]     OE_DATA_83_const_net_27;
wire   [3:0]     OE_DATA_84_const_net_27;
wire   [3:0]     OE_DATA_85_const_net_27;
wire   [3:0]     OE_DATA_86_const_net_27;
wire   [3:0]     OE_DATA_87_const_net_27;
wire   [3:0]     OE_DATA_88_const_net_27;
wire   [3:0]     OE_DATA_89_const_net_27;
wire   [3:0]     OE_DATA_90_const_net_27;
wire   [3:0]     OE_DATA_91_const_net_27;
wire   [3:0]     OE_DATA_92_const_net_27;
wire   [3:0]     OE_DATA_93_const_net_27;
wire   [3:0]     OE_DATA_94_const_net_27;
wire   [3:0]     OE_DATA_95_const_net_27;
wire   [3:0]     OE_DATA_96_const_net_27;
wire   [3:0]     OE_DATA_97_const_net_27;
wire   [3:0]     OE_DATA_98_const_net_27;
wire   [3:0]     OE_DATA_99_const_net_27;
wire   [3:0]     OE_DATA_100_const_net_27;
wire   [3:0]     OE_DATA_101_const_net_27;
wire   [3:0]     OE_DATA_102_const_net_27;
wire   [3:0]     OE_DATA_103_const_net_27;
wire   [3:0]     OE_DATA_104_const_net_27;
wire   [3:0]     OE_DATA_105_const_net_27;
wire   [3:0]     OE_DATA_106_const_net_27;
wire   [3:0]     OE_DATA_107_const_net_27;
wire   [3:0]     OE_DATA_108_const_net_27;
wire   [3:0]     OE_DATA_109_const_net_27;
wire   [3:0]     OE_DATA_110_const_net_27;
wire   [3:0]     OE_DATA_111_const_net_27;
wire   [3:0]     OE_DATA_112_const_net_27;
wire   [3:0]     OE_DATA_113_const_net_27;
wire   [3:0]     OE_DATA_114_const_net_27;
wire   [3:0]     OE_DATA_115_const_net_27;
wire   [3:0]     OE_DATA_116_const_net_27;
wire   [3:0]     OE_DATA_117_const_net_27;
wire   [3:0]     OE_DATA_118_const_net_27;
wire   [3:0]     OE_DATA_119_const_net_27;
wire   [3:0]     OE_DATA_120_const_net_27;
wire   [3:0]     OE_DATA_121_const_net_27;
wire   [3:0]     OE_DATA_122_const_net_27;
wire   [3:0]     OE_DATA_123_const_net_27;
wire   [3:0]     OE_DATA_124_const_net_27;
wire   [3:0]     OE_DATA_125_const_net_27;
wire   [3:0]     OE_DATA_126_const_net_27;
wire   [3:0]     OE_DATA_127_const_net_27;
wire   [1:0]     RX_DQS_90_const_net_19;
wire   [2:0]     FIFO_WR_PTR_const_net_20;
wire   [2:0]     FIFO_RD_PTR_const_net_20;
wire   [2:0]     EYE_MONITOR_LANE_WIDTH_const_net_22;
wire   [1:0]     TX_DATA_1_const_net_22;
wire   [1:0]     TX_DATA_2_const_net_24;
wire   [1:0]     TX_DATA_3_const_net_24;
wire   [1:0]     TX_DATA_4_const_net_24;
wire   [1:0]     TX_DATA_5_const_net_24;
wire   [1:0]     TX_DATA_6_const_net_24;
wire   [1:0]     TX_DATA_7_const_net_24;
wire   [1:0]     TX_DATA_8_const_net_27;
wire   [1:0]     TX_DATA_9_const_net_27;
wire   [1:0]     TX_DATA_10_const_net_27;
wire   [1:0]     TX_DATA_11_const_net_27;
wire   [1:0]     TX_DATA_12_const_net_28;
wire   [1:0]     TX_DATA_13_const_net_28;
wire   [1:0]     TX_DATA_14_const_net_28;
wire   [1:0]     TX_DATA_15_const_net_28;
wire   [1:0]     TX_DATA_16_const_net_28;
wire   [1:0]     TX_DATA_17_const_net_28;
wire   [1:0]     TX_DATA_18_const_net_28;
wire   [1:0]     TX_DATA_19_const_net_28;
wire   [1:0]     TX_DATA_20_const_net_28;
wire   [1:0]     TX_DATA_21_const_net_28;
wire   [1:0]     TX_DATA_22_const_net_28;
wire   [1:0]     TX_DATA_23_const_net_28;
wire   [1:0]     TX_DATA_24_const_net_28;
wire   [1:0]     TX_DATA_25_const_net_28;
wire   [1:0]     TX_DATA_26_const_net_28;
wire   [1:0]     TX_DATA_27_const_net_28;
wire   [1:0]     TX_DATA_28_const_net_28;
wire   [1:0]     TX_DATA_29_const_net_28;
wire   [1:0]     TX_DATA_30_const_net_28;
wire   [1:0]     TX_DATA_31_const_net_28;
wire   [1:0]     TX_DATA_32_const_net_28;
wire   [1:0]     TX_DATA_33_const_net_28;
wire   [1:0]     TX_DATA_34_const_net_28;
wire   [1:0]     TX_DATA_35_const_net_28;
wire   [1:0]     TX_DATA_36_const_net_28;
wire   [1:0]     TX_DATA_37_const_net_28;
wire   [1:0]     TX_DATA_38_const_net_28;
wire   [1:0]     TX_DATA_39_const_net_28;
wire   [1:0]     TX_DATA_40_const_net_28;
wire   [1:0]     TX_DATA_41_const_net_28;
wire   [1:0]     TX_DATA_42_const_net_28;
wire   [1:0]     TX_DATA_43_const_net_28;
wire   [1:0]     TX_DATA_44_const_net_28;
wire   [1:0]     TX_DATA_45_const_net_28;
wire   [1:0]     TX_DATA_46_const_net_28;
wire   [1:0]     TX_DATA_47_const_net_28;
wire   [1:0]     TX_DATA_48_const_net_28;
wire   [1:0]     TX_DATA_49_const_net_28;
wire   [1:0]     TX_DATA_50_const_net_28;
wire   [1:0]     TX_DATA_51_const_net_28;
wire   [1:0]     TX_DATA_52_const_net_28;
wire   [1:0]     TX_DATA_53_const_net_28;
wire   [1:0]     TX_DATA_54_const_net_28;
wire   [1:0]     TX_DATA_55_const_net_28;
wire   [1:0]     TX_DATA_56_const_net_28;
wire   [1:0]     TX_DATA_57_const_net_28;
wire   [1:0]     TX_DATA_58_const_net_28;
wire   [1:0]     TX_DATA_59_const_net_28;
wire   [1:0]     TX_DATA_60_const_net_28;
wire   [1:0]     TX_DATA_61_const_net_28;
wire   [1:0]     TX_DATA_62_const_net_28;
wire   [1:0]     TX_DATA_63_const_net_28;
wire   [1:0]     TX_DATA_64_const_net_28;
wire   [1:0]     TX_DATA_65_const_net_28;
wire   [1:0]     TX_DATA_66_const_net_28;
wire   [1:0]     TX_DATA_67_const_net_28;
wire   [1:0]     TX_DATA_68_const_net_28;
wire   [1:0]     TX_DATA_69_const_net_28;
wire   [1:0]     TX_DATA_70_const_net_28;
wire   [1:0]     TX_DATA_71_const_net_28;
wire   [1:0]     TX_DATA_72_const_net_28;
wire   [1:0]     TX_DATA_73_const_net_28;
wire   [1:0]     TX_DATA_74_const_net_28;
wire   [1:0]     TX_DATA_75_const_net_28;
wire   [1:0]     TX_DATA_76_const_net_28;
wire   [1:0]     TX_DATA_77_const_net_28;
wire   [1:0]     TX_DATA_78_const_net_28;
wire   [1:0]     TX_DATA_79_const_net_28;
wire   [1:0]     TX_DATA_80_const_net_28;
wire   [1:0]     TX_DATA_81_const_net_28;
wire   [1:0]     TX_DATA_82_const_net_28;
wire   [1:0]     TX_DATA_83_const_net_28;
wire   [1:0]     TX_DATA_84_const_net_28;
wire   [1:0]     TX_DATA_85_const_net_28;
wire   [1:0]     TX_DATA_86_const_net_28;
wire   [1:0]     TX_DATA_87_const_net_28;
wire   [1:0]     TX_DATA_88_const_net_28;
wire   [1:0]     TX_DATA_89_const_net_28;
wire   [1:0]     TX_DATA_90_const_net_28;
wire   [1:0]     TX_DATA_91_const_net_28;
wire   [1:0]     TX_DATA_92_const_net_28;
wire   [1:0]     TX_DATA_93_const_net_28;
wire   [1:0]     TX_DATA_94_const_net_28;
wire   [1:0]     TX_DATA_95_const_net_28;
wire   [1:0]     TX_DATA_96_const_net_28;
wire   [1:0]     TX_DATA_97_const_net_28;
wire   [1:0]     TX_DATA_98_const_net_28;
wire   [1:0]     TX_DATA_99_const_net_28;
wire   [1:0]     TX_DATA_100_const_net_28;
wire   [1:0]     TX_DATA_101_const_net_28;
wire   [1:0]     TX_DATA_102_const_net_28;
wire   [1:0]     TX_DATA_103_const_net_28;
wire   [1:0]     TX_DATA_104_const_net_28;
wire   [1:0]     TX_DATA_105_const_net_28;
wire   [1:0]     TX_DATA_106_const_net_28;
wire   [1:0]     TX_DATA_107_const_net_28;
wire   [1:0]     TX_DATA_108_const_net_28;
wire   [1:0]     TX_DATA_109_const_net_28;
wire   [1:0]     TX_DATA_110_const_net_28;
wire   [1:0]     TX_DATA_111_const_net_28;
wire   [1:0]     TX_DATA_112_const_net_28;
wire   [1:0]     TX_DATA_113_const_net_28;
wire   [1:0]     TX_DATA_114_const_net_28;
wire   [1:0]     TX_DATA_115_const_net_28;
wire   [1:0]     TX_DATA_116_const_net_28;
wire   [1:0]     TX_DATA_117_const_net_28;
wire   [1:0]     TX_DATA_118_const_net_28;
wire   [1:0]     TX_DATA_119_const_net_28;
wire   [1:0]     TX_DATA_120_const_net_28;
wire   [1:0]     TX_DATA_121_const_net_28;
wire   [1:0]     TX_DATA_122_const_net_28;
wire   [1:0]     TX_DATA_123_const_net_28;
wire   [1:0]     TX_DATA_124_const_net_28;
wire   [1:0]     TX_DATA_125_const_net_28;
wire   [1:0]     TX_DATA_126_const_net_28;
wire   [1:0]     TX_DATA_127_const_net_28;
wire   [1:0]     OE_DATA_1_const_net_25;
wire   [1:0]     OE_DATA_2_const_net_25;
wire   [1:0]     OE_DATA_3_const_net_25;
wire   [1:0]     OE_DATA_4_const_net_25;
wire   [1:0]     OE_DATA_5_const_net_25;
wire   [1:0]     OE_DATA_6_const_net_25;
wire   [1:0]     OE_DATA_7_const_net_25;
wire   [1:0]     OE_DATA_8_const_net_28;
wire   [1:0]     OE_DATA_9_const_net_28;
wire   [1:0]     OE_DATA_10_const_net_28;
wire   [1:0]     OE_DATA_11_const_net_28;
wire   [1:0]     OE_DATA_12_const_net_28;
wire   [1:0]     OE_DATA_13_const_net_28;
wire   [1:0]     OE_DATA_14_const_net_28;
wire   [1:0]     OE_DATA_15_const_net_28;
wire   [1:0]     OE_DATA_16_const_net_28;
wire   [1:0]     OE_DATA_17_const_net_28;
wire   [1:0]     OE_DATA_18_const_net_28;
wire   [1:0]     OE_DATA_19_const_net_28;
wire   [1:0]     OE_DATA_20_const_net_28;
wire   [1:0]     OE_DATA_21_const_net_28;
wire   [1:0]     OE_DATA_22_const_net_28;
wire   [1:0]     OE_DATA_23_const_net_28;
wire   [1:0]     OE_DATA_24_const_net_28;
wire   [1:0]     OE_DATA_25_const_net_28;
wire   [1:0]     OE_DATA_26_const_net_28;
wire   [1:0]     OE_DATA_27_const_net_28;
wire   [1:0]     OE_DATA_28_const_net_28;
wire   [1:0]     OE_DATA_29_const_net_28;
wire   [1:0]     OE_DATA_30_const_net_28;
wire   [1:0]     OE_DATA_31_const_net_28;
wire   [1:0]     OE_DATA_32_const_net_28;
wire   [1:0]     OE_DATA_33_const_net_28;
wire   [1:0]     OE_DATA_34_const_net_28;
wire   [1:0]     OE_DATA_35_const_net_28;
wire   [1:0]     OE_DATA_36_const_net_28;
wire   [1:0]     OE_DATA_37_const_net_28;
wire   [1:0]     OE_DATA_38_const_net_28;
wire   [1:0]     OE_DATA_39_const_net_28;
wire   [1:0]     OE_DATA_40_const_net_28;
wire   [1:0]     OE_DATA_41_const_net_28;
wire   [1:0]     OE_DATA_42_const_net_28;
wire   [1:0]     OE_DATA_43_const_net_28;
wire   [1:0]     OE_DATA_44_const_net_28;
wire   [1:0]     OE_DATA_45_const_net_28;
wire   [1:0]     OE_DATA_46_const_net_28;
wire   [1:0]     OE_DATA_47_const_net_28;
wire   [1:0]     OE_DATA_48_const_net_28;
wire   [1:0]     OE_DATA_49_const_net_28;
wire   [1:0]     OE_DATA_50_const_net_28;
wire   [1:0]     OE_DATA_51_const_net_28;
wire   [1:0]     OE_DATA_52_const_net_28;
wire   [1:0]     OE_DATA_53_const_net_28;
wire   [1:0]     OE_DATA_54_const_net_28;
wire   [1:0]     OE_DATA_55_const_net_28;
wire   [1:0]     OE_DATA_56_const_net_28;
wire   [1:0]     OE_DATA_57_const_net_28;
wire   [1:0]     OE_DATA_58_const_net_28;
wire   [1:0]     OE_DATA_59_const_net_28;
wire   [1:0]     OE_DATA_60_const_net_28;
wire   [1:0]     OE_DATA_61_const_net_28;
wire   [1:0]     OE_DATA_62_const_net_28;
wire   [1:0]     OE_DATA_63_const_net_28;
wire   [1:0]     OE_DATA_64_const_net_28;
wire   [1:0]     OE_DATA_65_const_net_28;
wire   [1:0]     OE_DATA_66_const_net_28;
wire   [1:0]     OE_DATA_67_const_net_28;
wire   [1:0]     OE_DATA_68_const_net_28;
wire   [1:0]     OE_DATA_69_const_net_28;
wire   [1:0]     OE_DATA_70_const_net_28;
wire   [1:0]     OE_DATA_71_const_net_28;
wire   [1:0]     OE_DATA_72_const_net_28;
wire   [1:0]     OE_DATA_73_const_net_28;
wire   [1:0]     OE_DATA_74_const_net_28;
wire   [1:0]     OE_DATA_75_const_net_28;
wire   [1:0]     OE_DATA_76_const_net_28;
wire   [1:0]     OE_DATA_77_const_net_28;
wire   [1:0]     OE_DATA_78_const_net_28;
wire   [1:0]     OE_DATA_79_const_net_28;
wire   [1:0]     OE_DATA_80_const_net_28;
wire   [1:0]     OE_DATA_81_const_net_28;
wire   [1:0]     OE_DATA_82_const_net_28;
wire   [1:0]     OE_DATA_83_const_net_28;
wire   [1:0]     OE_DATA_84_const_net_28;
wire   [1:0]     OE_DATA_85_const_net_28;
wire   [1:0]     OE_DATA_86_const_net_28;
wire   [1:0]     OE_DATA_87_const_net_28;
wire   [1:0]     OE_DATA_88_const_net_28;
wire   [1:0]     OE_DATA_89_const_net_28;
wire   [1:0]     OE_DATA_90_const_net_28;
wire   [1:0]     OE_DATA_91_const_net_28;
wire   [1:0]     OE_DATA_92_const_net_28;
wire   [1:0]     OE_DATA_93_const_net_28;
wire   [1:0]     OE_DATA_94_const_net_28;
wire   [1:0]     OE_DATA_95_const_net_28;
wire   [1:0]     OE_DATA_96_const_net_28;
wire   [1:0]     OE_DATA_97_const_net_28;
wire   [1:0]     OE_DATA_98_const_net_28;
wire   [1:0]     OE_DATA_99_const_net_28;
wire   [1:0]     OE_DATA_100_const_net_28;
wire   [1:0]     OE_DATA_101_const_net_28;
wire   [1:0]     OE_DATA_102_const_net_28;
wire   [1:0]     OE_DATA_103_const_net_28;
wire   [1:0]     OE_DATA_104_const_net_28;
wire   [1:0]     OE_DATA_105_const_net_28;
wire   [1:0]     OE_DATA_106_const_net_28;
wire   [1:0]     OE_DATA_107_const_net_28;
wire   [1:0]     OE_DATA_108_const_net_28;
wire   [1:0]     OE_DATA_109_const_net_28;
wire   [1:0]     OE_DATA_110_const_net_28;
wire   [1:0]     OE_DATA_111_const_net_28;
wire   [1:0]     OE_DATA_112_const_net_28;
wire   [1:0]     OE_DATA_113_const_net_28;
wire   [1:0]     OE_DATA_114_const_net_28;
wire   [1:0]     OE_DATA_115_const_net_28;
wire   [1:0]     OE_DATA_116_const_net_28;
wire   [1:0]     OE_DATA_117_const_net_28;
wire   [1:0]     OE_DATA_118_const_net_28;
wire   [1:0]     OE_DATA_119_const_net_28;
wire   [1:0]     OE_DATA_120_const_net_28;
wire   [1:0]     OE_DATA_121_const_net_28;
wire   [1:0]     OE_DATA_122_const_net_28;
wire   [1:0]     OE_DATA_123_const_net_28;
wire   [1:0]     OE_DATA_124_const_net_28;
wire   [1:0]     OE_DATA_125_const_net_28;
wire   [1:0]     OE_DATA_126_const_net_28;
wire   [1:0]     OE_DATA_127_const_net_28;
wire   [1:0]     RX_DQS_90_const_net_20;
wire   [2:0]     EYE_MONITOR_LANE_WIDTH_const_net_23;
wire   [7:0]     TX_DATA_1_const_net_23;
wire   [7:0]     TX_DATA_2_const_net_25;
wire   [7:0]     TX_DATA_3_const_net_25;
wire   [7:0]     TX_DATA_4_const_net_25;
wire   [7:0]     TX_DATA_5_const_net_25;
wire   [7:0]     TX_DATA_6_const_net_25;
wire   [7:0]     TX_DATA_7_const_net_25;
wire   [7:0]     TX_DATA_8_const_net_28;
wire   [7:0]     TX_DATA_9_const_net_28;
wire   [7:0]     TX_DATA_10_const_net_28;
wire   [7:0]     TX_DATA_11_const_net_28;
wire   [7:0]     TX_DATA_12_const_net_29;
wire   [7:0]     TX_DATA_13_const_net_29;
wire   [7:0]     TX_DATA_14_const_net_29;
wire   [7:0]     TX_DATA_15_const_net_29;
wire   [7:0]     TX_DATA_16_const_net_29;
wire   [7:0]     TX_DATA_17_const_net_29;
wire   [7:0]     TX_DATA_18_const_net_29;
wire   [7:0]     TX_DATA_19_const_net_29;
wire   [7:0]     TX_DATA_20_const_net_29;
wire   [7:0]     TX_DATA_21_const_net_29;
wire   [7:0]     TX_DATA_22_const_net_29;
wire   [7:0]     TX_DATA_23_const_net_29;
wire   [7:0]     TX_DATA_24_const_net_29;
wire   [7:0]     TX_DATA_25_const_net_29;
wire   [7:0]     TX_DATA_26_const_net_29;
wire   [7:0]     TX_DATA_27_const_net_29;
wire   [7:0]     TX_DATA_28_const_net_29;
wire   [7:0]     TX_DATA_29_const_net_29;
wire   [7:0]     TX_DATA_30_const_net_29;
wire   [7:0]     TX_DATA_31_const_net_29;
wire   [7:0]     TX_DATA_32_const_net_29;
wire   [7:0]     TX_DATA_33_const_net_29;
wire   [7:0]     TX_DATA_34_const_net_29;
wire   [7:0]     TX_DATA_35_const_net_29;
wire   [7:0]     TX_DATA_36_const_net_29;
wire   [7:0]     TX_DATA_37_const_net_29;
wire   [7:0]     TX_DATA_38_const_net_29;
wire   [7:0]     TX_DATA_39_const_net_29;
wire   [7:0]     TX_DATA_40_const_net_29;
wire   [7:0]     TX_DATA_41_const_net_29;
wire   [7:0]     TX_DATA_42_const_net_29;
wire   [7:0]     TX_DATA_43_const_net_29;
wire   [7:0]     TX_DATA_44_const_net_29;
wire   [7:0]     TX_DATA_45_const_net_29;
wire   [7:0]     TX_DATA_46_const_net_29;
wire   [7:0]     TX_DATA_47_const_net_29;
wire   [7:0]     TX_DATA_48_const_net_29;
wire   [7:0]     TX_DATA_49_const_net_29;
wire   [7:0]     TX_DATA_50_const_net_29;
wire   [7:0]     TX_DATA_51_const_net_29;
wire   [7:0]     TX_DATA_52_const_net_29;
wire   [7:0]     TX_DATA_53_const_net_29;
wire   [7:0]     TX_DATA_54_const_net_29;
wire   [7:0]     TX_DATA_55_const_net_29;
wire   [7:0]     TX_DATA_56_const_net_29;
wire   [7:0]     TX_DATA_57_const_net_29;
wire   [7:0]     TX_DATA_58_const_net_29;
wire   [7:0]     TX_DATA_59_const_net_29;
wire   [7:0]     TX_DATA_60_const_net_29;
wire   [7:0]     TX_DATA_61_const_net_29;
wire   [7:0]     TX_DATA_62_const_net_29;
wire   [7:0]     TX_DATA_63_const_net_29;
wire   [7:0]     TX_DATA_64_const_net_29;
wire   [7:0]     TX_DATA_65_const_net_29;
wire   [7:0]     TX_DATA_66_const_net_29;
wire   [7:0]     TX_DATA_67_const_net_29;
wire   [7:0]     TX_DATA_68_const_net_29;
wire   [7:0]     TX_DATA_69_const_net_29;
wire   [7:0]     TX_DATA_70_const_net_29;
wire   [7:0]     TX_DATA_71_const_net_29;
wire   [7:0]     TX_DATA_72_const_net_29;
wire   [7:0]     TX_DATA_73_const_net_29;
wire   [7:0]     TX_DATA_74_const_net_29;
wire   [7:0]     TX_DATA_75_const_net_29;
wire   [7:0]     TX_DATA_76_const_net_29;
wire   [7:0]     TX_DATA_77_const_net_29;
wire   [7:0]     TX_DATA_78_const_net_29;
wire   [7:0]     TX_DATA_79_const_net_29;
wire   [7:0]     TX_DATA_80_const_net_29;
wire   [7:0]     TX_DATA_81_const_net_29;
wire   [7:0]     TX_DATA_82_const_net_29;
wire   [7:0]     TX_DATA_83_const_net_29;
wire   [7:0]     TX_DATA_84_const_net_29;
wire   [7:0]     TX_DATA_85_const_net_29;
wire   [7:0]     TX_DATA_86_const_net_29;
wire   [7:0]     TX_DATA_87_const_net_29;
wire   [7:0]     TX_DATA_88_const_net_29;
wire   [7:0]     TX_DATA_89_const_net_29;
wire   [7:0]     TX_DATA_90_const_net_29;
wire   [7:0]     TX_DATA_91_const_net_29;
wire   [7:0]     TX_DATA_92_const_net_29;
wire   [7:0]     TX_DATA_93_const_net_29;
wire   [7:0]     TX_DATA_94_const_net_29;
wire   [7:0]     TX_DATA_95_const_net_29;
wire   [7:0]     TX_DATA_96_const_net_29;
wire   [7:0]     TX_DATA_97_const_net_29;
wire   [7:0]     TX_DATA_98_const_net_29;
wire   [7:0]     TX_DATA_99_const_net_29;
wire   [7:0]     TX_DATA_100_const_net_29;
wire   [7:0]     TX_DATA_101_const_net_29;
wire   [7:0]     TX_DATA_102_const_net_29;
wire   [7:0]     TX_DATA_103_const_net_29;
wire   [7:0]     TX_DATA_104_const_net_29;
wire   [7:0]     TX_DATA_105_const_net_29;
wire   [7:0]     TX_DATA_106_const_net_29;
wire   [7:0]     TX_DATA_107_const_net_29;
wire   [7:0]     TX_DATA_108_const_net_29;
wire   [7:0]     TX_DATA_109_const_net_29;
wire   [7:0]     TX_DATA_110_const_net_29;
wire   [7:0]     TX_DATA_111_const_net_29;
wire   [7:0]     TX_DATA_112_const_net_29;
wire   [7:0]     TX_DATA_113_const_net_29;
wire   [7:0]     TX_DATA_114_const_net_29;
wire   [7:0]     TX_DATA_115_const_net_29;
wire   [7:0]     TX_DATA_116_const_net_29;
wire   [7:0]     TX_DATA_117_const_net_29;
wire   [7:0]     TX_DATA_118_const_net_29;
wire   [7:0]     TX_DATA_119_const_net_29;
wire   [7:0]     TX_DATA_120_const_net_29;
wire   [7:0]     TX_DATA_121_const_net_29;
wire   [7:0]     TX_DATA_122_const_net_29;
wire   [7:0]     TX_DATA_123_const_net_29;
wire   [7:0]     TX_DATA_124_const_net_29;
wire   [7:0]     TX_DATA_125_const_net_29;
wire   [7:0]     TX_DATA_126_const_net_29;
wire   [7:0]     TX_DATA_127_const_net_29;
wire   [3:0]     OE_DATA_1_const_net_26;
wire   [3:0]     OE_DATA_2_const_net_26;
wire   [3:0]     OE_DATA_3_const_net_26;
wire   [3:0]     OE_DATA_4_const_net_26;
wire   [3:0]     OE_DATA_5_const_net_26;
wire   [3:0]     OE_DATA_6_const_net_26;
wire   [3:0]     OE_DATA_7_const_net_26;
wire   [3:0]     OE_DATA_8_const_net_29;
wire   [3:0]     OE_DATA_9_const_net_29;
wire   [3:0]     OE_DATA_10_const_net_29;
wire   [3:0]     OE_DATA_11_const_net_29;
wire   [3:0]     OE_DATA_12_const_net_29;
wire   [3:0]     OE_DATA_13_const_net_29;
wire   [3:0]     OE_DATA_14_const_net_29;
wire   [3:0]     OE_DATA_15_const_net_29;
wire   [3:0]     OE_DATA_16_const_net_29;
wire   [3:0]     OE_DATA_17_const_net_29;
wire   [3:0]     OE_DATA_18_const_net_29;
wire   [3:0]     OE_DATA_19_const_net_29;
wire   [3:0]     OE_DATA_20_const_net_29;
wire   [3:0]     OE_DATA_21_const_net_29;
wire   [3:0]     OE_DATA_22_const_net_29;
wire   [3:0]     OE_DATA_23_const_net_29;
wire   [3:0]     OE_DATA_24_const_net_29;
wire   [3:0]     OE_DATA_25_const_net_29;
wire   [3:0]     OE_DATA_26_const_net_29;
wire   [3:0]     OE_DATA_27_const_net_29;
wire   [3:0]     OE_DATA_28_const_net_29;
wire   [3:0]     OE_DATA_29_const_net_29;
wire   [3:0]     OE_DATA_30_const_net_29;
wire   [3:0]     OE_DATA_31_const_net_29;
wire   [3:0]     OE_DATA_32_const_net_29;
wire   [3:0]     OE_DATA_33_const_net_29;
wire   [3:0]     OE_DATA_34_const_net_29;
wire   [3:0]     OE_DATA_35_const_net_29;
wire   [3:0]     OE_DATA_36_const_net_29;
wire   [3:0]     OE_DATA_37_const_net_29;
wire   [3:0]     OE_DATA_38_const_net_29;
wire   [3:0]     OE_DATA_39_const_net_29;
wire   [3:0]     OE_DATA_40_const_net_29;
wire   [3:0]     OE_DATA_41_const_net_29;
wire   [3:0]     OE_DATA_42_const_net_29;
wire   [3:0]     OE_DATA_43_const_net_29;
wire   [3:0]     OE_DATA_44_const_net_29;
wire   [3:0]     OE_DATA_45_const_net_29;
wire   [3:0]     OE_DATA_46_const_net_29;
wire   [3:0]     OE_DATA_47_const_net_29;
wire   [3:0]     OE_DATA_48_const_net_29;
wire   [3:0]     OE_DATA_49_const_net_29;
wire   [3:0]     OE_DATA_50_const_net_29;
wire   [3:0]     OE_DATA_51_const_net_29;
wire   [3:0]     OE_DATA_52_const_net_29;
wire   [3:0]     OE_DATA_53_const_net_29;
wire   [3:0]     OE_DATA_54_const_net_29;
wire   [3:0]     OE_DATA_55_const_net_29;
wire   [3:0]     OE_DATA_56_const_net_29;
wire   [3:0]     OE_DATA_57_const_net_29;
wire   [3:0]     OE_DATA_58_const_net_29;
wire   [3:0]     OE_DATA_59_const_net_29;
wire   [3:0]     OE_DATA_60_const_net_29;
wire   [3:0]     OE_DATA_61_const_net_29;
wire   [3:0]     OE_DATA_62_const_net_29;
wire   [3:0]     OE_DATA_63_const_net_29;
wire   [3:0]     OE_DATA_64_const_net_29;
wire   [3:0]     OE_DATA_65_const_net_29;
wire   [3:0]     OE_DATA_66_const_net_29;
wire   [3:0]     OE_DATA_67_const_net_29;
wire   [3:0]     OE_DATA_68_const_net_29;
wire   [3:0]     OE_DATA_69_const_net_29;
wire   [3:0]     OE_DATA_70_const_net_29;
wire   [3:0]     OE_DATA_71_const_net_29;
wire   [3:0]     OE_DATA_72_const_net_29;
wire   [3:0]     OE_DATA_73_const_net_29;
wire   [3:0]     OE_DATA_74_const_net_29;
wire   [3:0]     OE_DATA_75_const_net_29;
wire   [3:0]     OE_DATA_76_const_net_29;
wire   [3:0]     OE_DATA_77_const_net_29;
wire   [3:0]     OE_DATA_78_const_net_29;
wire   [3:0]     OE_DATA_79_const_net_29;
wire   [3:0]     OE_DATA_80_const_net_29;
wire   [3:0]     OE_DATA_81_const_net_29;
wire   [3:0]     OE_DATA_82_const_net_29;
wire   [3:0]     OE_DATA_83_const_net_29;
wire   [3:0]     OE_DATA_84_const_net_29;
wire   [3:0]     OE_DATA_85_const_net_29;
wire   [3:0]     OE_DATA_86_const_net_29;
wire   [3:0]     OE_DATA_87_const_net_29;
wire   [3:0]     OE_DATA_88_const_net_29;
wire   [3:0]     OE_DATA_89_const_net_29;
wire   [3:0]     OE_DATA_90_const_net_29;
wire   [3:0]     OE_DATA_91_const_net_29;
wire   [3:0]     OE_DATA_92_const_net_29;
wire   [3:0]     OE_DATA_93_const_net_29;
wire   [3:0]     OE_DATA_94_const_net_29;
wire   [3:0]     OE_DATA_95_const_net_29;
wire   [3:0]     OE_DATA_96_const_net_29;
wire   [3:0]     OE_DATA_97_const_net_29;
wire   [3:0]     OE_DATA_98_const_net_29;
wire   [3:0]     OE_DATA_99_const_net_29;
wire   [3:0]     OE_DATA_100_const_net_29;
wire   [3:0]     OE_DATA_101_const_net_29;
wire   [3:0]     OE_DATA_102_const_net_29;
wire   [3:0]     OE_DATA_103_const_net_29;
wire   [3:0]     OE_DATA_104_const_net_29;
wire   [3:0]     OE_DATA_105_const_net_29;
wire   [3:0]     OE_DATA_106_const_net_29;
wire   [3:0]     OE_DATA_107_const_net_29;
wire   [3:0]     OE_DATA_108_const_net_29;
wire   [3:0]     OE_DATA_109_const_net_29;
wire   [3:0]     OE_DATA_110_const_net_29;
wire   [3:0]     OE_DATA_111_const_net_29;
wire   [3:0]     OE_DATA_112_const_net_29;
wire   [3:0]     OE_DATA_113_const_net_29;
wire   [3:0]     OE_DATA_114_const_net_29;
wire   [3:0]     OE_DATA_115_const_net_29;
wire   [3:0]     OE_DATA_116_const_net_29;
wire   [3:0]     OE_DATA_117_const_net_29;
wire   [3:0]     OE_DATA_118_const_net_29;
wire   [3:0]     OE_DATA_119_const_net_29;
wire   [3:0]     OE_DATA_120_const_net_29;
wire   [3:0]     OE_DATA_121_const_net_29;
wire   [3:0]     OE_DATA_122_const_net_29;
wire   [3:0]     OE_DATA_123_const_net_29;
wire   [3:0]     OE_DATA_124_const_net_29;
wire   [3:0]     OE_DATA_125_const_net_29;
wire   [3:0]     OE_DATA_126_const_net_29;
wire   [3:0]     OE_DATA_127_const_net_29;
wire   [10:0]    CDR_CLK_B_SEL_const_net_3;
wire   [2:0]     FIFO_WR_PTR_const_net_21;
wire   [2:0]     FIFO_RD_PTR_const_net_21;
wire   [2:0]     EYE_MONITOR_LANE_WIDTH_const_net_24;
wire   [7:0]     TX_DATA_1_const_net_24;
wire   [7:0]     TX_DATA_2_const_net_26;
wire   [7:0]     TX_DATA_3_const_net_26;
wire   [7:0]     TX_DATA_4_const_net_26;
wire   [7:0]     TX_DATA_5_const_net_26;
wire   [7:0]     TX_DATA_6_const_net_26;
wire   [7:0]     TX_DATA_7_const_net_26;
wire   [7:0]     TX_DATA_8_const_net_29;
wire   [7:0]     TX_DATA_9_const_net_29;
wire   [7:0]     TX_DATA_10_const_net_29;
wire   [7:0]     TX_DATA_11_const_net_29;
wire   [7:0]     TX_DATA_12_const_net_30;
wire   [7:0]     TX_DATA_13_const_net_30;
wire   [7:0]     TX_DATA_14_const_net_30;
wire   [7:0]     TX_DATA_15_const_net_30;
wire   [7:0]     TX_DATA_16_const_net_30;
wire   [7:0]     TX_DATA_17_const_net_30;
wire   [7:0]     TX_DATA_18_const_net_30;
wire   [7:0]     TX_DATA_19_const_net_30;
wire   [7:0]     TX_DATA_20_const_net_30;
wire   [7:0]     TX_DATA_21_const_net_30;
wire   [7:0]     TX_DATA_22_const_net_30;
wire   [7:0]     TX_DATA_23_const_net_30;
wire   [7:0]     TX_DATA_24_const_net_30;
wire   [7:0]     TX_DATA_25_const_net_30;
wire   [7:0]     TX_DATA_26_const_net_30;
wire   [7:0]     TX_DATA_27_const_net_30;
wire   [7:0]     TX_DATA_28_const_net_30;
wire   [7:0]     TX_DATA_29_const_net_30;
wire   [7:0]     TX_DATA_30_const_net_30;
wire   [7:0]     TX_DATA_31_const_net_30;
wire   [7:0]     TX_DATA_32_const_net_30;
wire   [7:0]     TX_DATA_33_const_net_30;
wire   [7:0]     TX_DATA_34_const_net_30;
wire   [7:0]     TX_DATA_35_const_net_30;
wire   [7:0]     TX_DATA_36_const_net_30;
wire   [7:0]     TX_DATA_37_const_net_30;
wire   [7:0]     TX_DATA_38_const_net_30;
wire   [7:0]     TX_DATA_39_const_net_30;
wire   [7:0]     TX_DATA_40_const_net_30;
wire   [7:0]     TX_DATA_41_const_net_30;
wire   [7:0]     TX_DATA_42_const_net_30;
wire   [7:0]     TX_DATA_43_const_net_30;
wire   [7:0]     TX_DATA_44_const_net_30;
wire   [7:0]     TX_DATA_45_const_net_30;
wire   [7:0]     TX_DATA_46_const_net_30;
wire   [7:0]     TX_DATA_47_const_net_30;
wire   [7:0]     TX_DATA_48_const_net_30;
wire   [7:0]     TX_DATA_49_const_net_30;
wire   [7:0]     TX_DATA_50_const_net_30;
wire   [7:0]     TX_DATA_51_const_net_30;
wire   [7:0]     TX_DATA_52_const_net_30;
wire   [7:0]     TX_DATA_53_const_net_30;
wire   [7:0]     TX_DATA_54_const_net_30;
wire   [7:0]     TX_DATA_55_const_net_30;
wire   [7:0]     TX_DATA_56_const_net_30;
wire   [7:0]     TX_DATA_57_const_net_30;
wire   [7:0]     TX_DATA_58_const_net_30;
wire   [7:0]     TX_DATA_59_const_net_30;
wire   [7:0]     TX_DATA_60_const_net_30;
wire   [7:0]     TX_DATA_61_const_net_30;
wire   [7:0]     TX_DATA_62_const_net_30;
wire   [7:0]     TX_DATA_63_const_net_30;
wire   [7:0]     TX_DATA_64_const_net_30;
wire   [7:0]     TX_DATA_65_const_net_30;
wire   [7:0]     TX_DATA_66_const_net_30;
wire   [7:0]     TX_DATA_67_const_net_30;
wire   [7:0]     TX_DATA_68_const_net_30;
wire   [7:0]     TX_DATA_69_const_net_30;
wire   [7:0]     TX_DATA_70_const_net_30;
wire   [7:0]     TX_DATA_71_const_net_30;
wire   [7:0]     TX_DATA_72_const_net_30;
wire   [7:0]     TX_DATA_73_const_net_30;
wire   [7:0]     TX_DATA_74_const_net_30;
wire   [7:0]     TX_DATA_75_const_net_30;
wire   [7:0]     TX_DATA_76_const_net_30;
wire   [7:0]     TX_DATA_77_const_net_30;
wire   [7:0]     TX_DATA_78_const_net_30;
wire   [7:0]     TX_DATA_79_const_net_30;
wire   [7:0]     TX_DATA_80_const_net_30;
wire   [7:0]     TX_DATA_81_const_net_30;
wire   [7:0]     TX_DATA_82_const_net_30;
wire   [7:0]     TX_DATA_83_const_net_30;
wire   [7:0]     TX_DATA_84_const_net_30;
wire   [7:0]     TX_DATA_85_const_net_30;
wire   [7:0]     TX_DATA_86_const_net_30;
wire   [7:0]     TX_DATA_87_const_net_30;
wire   [7:0]     TX_DATA_88_const_net_30;
wire   [7:0]     TX_DATA_89_const_net_30;
wire   [7:0]     TX_DATA_90_const_net_30;
wire   [7:0]     TX_DATA_91_const_net_30;
wire   [7:0]     TX_DATA_92_const_net_30;
wire   [7:0]     TX_DATA_93_const_net_30;
wire   [7:0]     TX_DATA_94_const_net_30;
wire   [7:0]     TX_DATA_95_const_net_30;
wire   [7:0]     TX_DATA_96_const_net_30;
wire   [7:0]     TX_DATA_97_const_net_30;
wire   [7:0]     TX_DATA_98_const_net_30;
wire   [7:0]     TX_DATA_99_const_net_30;
wire   [7:0]     TX_DATA_100_const_net_30;
wire   [7:0]     TX_DATA_101_const_net_30;
wire   [7:0]     TX_DATA_102_const_net_30;
wire   [7:0]     TX_DATA_103_const_net_30;
wire   [7:0]     TX_DATA_104_const_net_30;
wire   [7:0]     TX_DATA_105_const_net_30;
wire   [7:0]     TX_DATA_106_const_net_30;
wire   [7:0]     TX_DATA_107_const_net_30;
wire   [7:0]     TX_DATA_108_const_net_30;
wire   [7:0]     TX_DATA_109_const_net_30;
wire   [7:0]     TX_DATA_110_const_net_30;
wire   [7:0]     TX_DATA_111_const_net_30;
wire   [7:0]     TX_DATA_112_const_net_30;
wire   [7:0]     TX_DATA_113_const_net_30;
wire   [7:0]     TX_DATA_114_const_net_30;
wire   [7:0]     TX_DATA_115_const_net_30;
wire   [7:0]     TX_DATA_116_const_net_30;
wire   [7:0]     TX_DATA_117_const_net_30;
wire   [7:0]     TX_DATA_118_const_net_30;
wire   [7:0]     TX_DATA_119_const_net_30;
wire   [7:0]     TX_DATA_120_const_net_30;
wire   [7:0]     TX_DATA_121_const_net_30;
wire   [7:0]     TX_DATA_122_const_net_30;
wire   [7:0]     TX_DATA_123_const_net_30;
wire   [7:0]     TX_DATA_124_const_net_30;
wire   [7:0]     TX_DATA_125_const_net_30;
wire   [7:0]     TX_DATA_126_const_net_30;
wire   [7:0]     TX_DATA_127_const_net_30;
wire   [3:0]     OE_DATA_1_const_net_27;
wire   [3:0]     OE_DATA_2_const_net_27;
wire   [3:0]     OE_DATA_3_const_net_27;
wire   [3:0]     OE_DATA_4_const_net_27;
wire   [3:0]     OE_DATA_5_const_net_27;
wire   [3:0]     OE_DATA_6_const_net_27;
wire   [3:0]     OE_DATA_7_const_net_27;
wire   [3:0]     OE_DATA_8_const_net_30;
wire   [3:0]     OE_DATA_9_const_net_30;
wire   [3:0]     OE_DATA_10_const_net_30;
wire   [3:0]     OE_DATA_11_const_net_30;
wire   [3:0]     OE_DATA_12_const_net_30;
wire   [3:0]     OE_DATA_13_const_net_30;
wire   [3:0]     OE_DATA_14_const_net_30;
wire   [3:0]     OE_DATA_15_const_net_30;
wire   [3:0]     OE_DATA_16_const_net_30;
wire   [3:0]     OE_DATA_17_const_net_30;
wire   [3:0]     OE_DATA_18_const_net_30;
wire   [3:0]     OE_DATA_19_const_net_30;
wire   [3:0]     OE_DATA_20_const_net_30;
wire   [3:0]     OE_DATA_21_const_net_30;
wire   [3:0]     OE_DATA_22_const_net_30;
wire   [3:0]     OE_DATA_23_const_net_30;
wire   [3:0]     OE_DATA_24_const_net_30;
wire   [3:0]     OE_DATA_25_const_net_30;
wire   [3:0]     OE_DATA_26_const_net_30;
wire   [3:0]     OE_DATA_27_const_net_30;
wire   [3:0]     OE_DATA_28_const_net_30;
wire   [3:0]     OE_DATA_29_const_net_30;
wire   [3:0]     OE_DATA_30_const_net_30;
wire   [3:0]     OE_DATA_31_const_net_30;
wire   [3:0]     OE_DATA_32_const_net_30;
wire   [3:0]     OE_DATA_33_const_net_30;
wire   [3:0]     OE_DATA_34_const_net_30;
wire   [3:0]     OE_DATA_35_const_net_30;
wire   [3:0]     OE_DATA_36_const_net_30;
wire   [3:0]     OE_DATA_37_const_net_30;
wire   [3:0]     OE_DATA_38_const_net_30;
wire   [3:0]     OE_DATA_39_const_net_30;
wire   [3:0]     OE_DATA_40_const_net_30;
wire   [3:0]     OE_DATA_41_const_net_30;
wire   [3:0]     OE_DATA_42_const_net_30;
wire   [3:0]     OE_DATA_43_const_net_30;
wire   [3:0]     OE_DATA_44_const_net_30;
wire   [3:0]     OE_DATA_45_const_net_30;
wire   [3:0]     OE_DATA_46_const_net_30;
wire   [3:0]     OE_DATA_47_const_net_30;
wire   [3:0]     OE_DATA_48_const_net_30;
wire   [3:0]     OE_DATA_49_const_net_30;
wire   [3:0]     OE_DATA_50_const_net_30;
wire   [3:0]     OE_DATA_51_const_net_30;
wire   [3:0]     OE_DATA_52_const_net_30;
wire   [3:0]     OE_DATA_53_const_net_30;
wire   [3:0]     OE_DATA_54_const_net_30;
wire   [3:0]     OE_DATA_55_const_net_30;
wire   [3:0]     OE_DATA_56_const_net_30;
wire   [3:0]     OE_DATA_57_const_net_30;
wire   [3:0]     OE_DATA_58_const_net_30;
wire   [3:0]     OE_DATA_59_const_net_30;
wire   [3:0]     OE_DATA_60_const_net_30;
wire   [3:0]     OE_DATA_61_const_net_30;
wire   [3:0]     OE_DATA_62_const_net_30;
wire   [3:0]     OE_DATA_63_const_net_30;
wire   [3:0]     OE_DATA_64_const_net_30;
wire   [3:0]     OE_DATA_65_const_net_30;
wire   [3:0]     OE_DATA_66_const_net_30;
wire   [3:0]     OE_DATA_67_const_net_30;
wire   [3:0]     OE_DATA_68_const_net_30;
wire   [3:0]     OE_DATA_69_const_net_30;
wire   [3:0]     OE_DATA_70_const_net_30;
wire   [3:0]     OE_DATA_71_const_net_30;
wire   [3:0]     OE_DATA_72_const_net_30;
wire   [3:0]     OE_DATA_73_const_net_30;
wire   [3:0]     OE_DATA_74_const_net_30;
wire   [3:0]     OE_DATA_75_const_net_30;
wire   [3:0]     OE_DATA_76_const_net_30;
wire   [3:0]     OE_DATA_77_const_net_30;
wire   [3:0]     OE_DATA_78_const_net_30;
wire   [3:0]     OE_DATA_79_const_net_30;
wire   [3:0]     OE_DATA_80_const_net_30;
wire   [3:0]     OE_DATA_81_const_net_30;
wire   [3:0]     OE_DATA_82_const_net_30;
wire   [3:0]     OE_DATA_83_const_net_30;
wire   [3:0]     OE_DATA_84_const_net_30;
wire   [3:0]     OE_DATA_85_const_net_30;
wire   [3:0]     OE_DATA_86_const_net_30;
wire   [3:0]     OE_DATA_87_const_net_30;
wire   [3:0]     OE_DATA_88_const_net_30;
wire   [3:0]     OE_DATA_89_const_net_30;
wire   [3:0]     OE_DATA_90_const_net_30;
wire   [3:0]     OE_DATA_91_const_net_30;
wire   [3:0]     OE_DATA_92_const_net_30;
wire   [3:0]     OE_DATA_93_const_net_30;
wire   [3:0]     OE_DATA_94_const_net_30;
wire   [3:0]     OE_DATA_95_const_net_30;
wire   [3:0]     OE_DATA_96_const_net_30;
wire   [3:0]     OE_DATA_97_const_net_30;
wire   [3:0]     OE_DATA_98_const_net_30;
wire   [3:0]     OE_DATA_99_const_net_30;
wire   [3:0]     OE_DATA_100_const_net_30;
wire   [3:0]     OE_DATA_101_const_net_30;
wire   [3:0]     OE_DATA_102_const_net_30;
wire   [3:0]     OE_DATA_103_const_net_30;
wire   [3:0]     OE_DATA_104_const_net_30;
wire   [3:0]     OE_DATA_105_const_net_30;
wire   [3:0]     OE_DATA_106_const_net_30;
wire   [3:0]     OE_DATA_107_const_net_30;
wire   [3:0]     OE_DATA_108_const_net_30;
wire   [3:0]     OE_DATA_109_const_net_30;
wire   [3:0]     OE_DATA_110_const_net_30;
wire   [3:0]     OE_DATA_111_const_net_30;
wire   [3:0]     OE_DATA_112_const_net_30;
wire   [3:0]     OE_DATA_113_const_net_30;
wire   [3:0]     OE_DATA_114_const_net_30;
wire   [3:0]     OE_DATA_115_const_net_30;
wire   [3:0]     OE_DATA_116_const_net_30;
wire   [3:0]     OE_DATA_117_const_net_30;
wire   [3:0]     OE_DATA_118_const_net_30;
wire   [3:0]     OE_DATA_119_const_net_30;
wire   [3:0]     OE_DATA_120_const_net_30;
wire   [3:0]     OE_DATA_121_const_net_30;
wire   [3:0]     OE_DATA_122_const_net_30;
wire   [3:0]     OE_DATA_123_const_net_30;
wire   [3:0]     OE_DATA_124_const_net_30;
wire   [3:0]     OE_DATA_125_const_net_30;
wire   [3:0]     OE_DATA_126_const_net_30;
wire   [3:0]     OE_DATA_127_const_net_30;
wire   [7:0]     TX_DATA_8_const_net_30;
wire   [7:0]     TX_DATA_9_const_net_30;
wire   [7:0]     TX_DATA_10_const_net_30;
wire   [7:0]     TX_DATA_11_const_net_30;
wire   [7:0]     TX_DATA_12_const_net_31;
wire   [7:0]     TX_DATA_13_const_net_31;
wire   [7:0]     TX_DATA_14_const_net_31;
wire   [7:0]     TX_DATA_15_const_net_31;
wire   [7:0]     TX_DATA_16_const_net_31;
wire   [7:0]     TX_DATA_17_const_net_31;
wire   [7:0]     TX_DATA_18_const_net_31;
wire   [7:0]     TX_DATA_19_const_net_31;
wire   [7:0]     TX_DATA_20_const_net_31;
wire   [7:0]     TX_DATA_21_const_net_31;
wire   [7:0]     TX_DATA_22_const_net_31;
wire   [7:0]     TX_DATA_23_const_net_31;
wire   [7:0]     TX_DATA_24_const_net_31;
wire   [7:0]     TX_DATA_25_const_net_31;
wire   [7:0]     TX_DATA_26_const_net_31;
wire   [7:0]     TX_DATA_27_const_net_31;
wire   [7:0]     TX_DATA_28_const_net_31;
wire   [7:0]     TX_DATA_29_const_net_31;
wire   [7:0]     TX_DATA_30_const_net_31;
wire   [7:0]     TX_DATA_31_const_net_31;
wire   [7:0]     TX_DATA_32_const_net_31;
wire   [7:0]     TX_DATA_33_const_net_31;
wire   [7:0]     TX_DATA_34_const_net_31;
wire   [7:0]     TX_DATA_35_const_net_31;
wire   [7:0]     TX_DATA_36_const_net_31;
wire   [7:0]     TX_DATA_37_const_net_31;
wire   [7:0]     TX_DATA_38_const_net_31;
wire   [7:0]     TX_DATA_39_const_net_31;
wire   [7:0]     TX_DATA_40_const_net_31;
wire   [7:0]     TX_DATA_41_const_net_31;
wire   [7:0]     TX_DATA_42_const_net_31;
wire   [7:0]     TX_DATA_43_const_net_31;
wire   [7:0]     TX_DATA_44_const_net_31;
wire   [7:0]     TX_DATA_45_const_net_31;
wire   [7:0]     TX_DATA_46_const_net_31;
wire   [7:0]     TX_DATA_47_const_net_31;
wire   [7:0]     TX_DATA_48_const_net_31;
wire   [7:0]     TX_DATA_49_const_net_31;
wire   [7:0]     TX_DATA_50_const_net_31;
wire   [7:0]     TX_DATA_51_const_net_31;
wire   [7:0]     TX_DATA_52_const_net_31;
wire   [7:0]     TX_DATA_53_const_net_31;
wire   [7:0]     TX_DATA_54_const_net_31;
wire   [7:0]     TX_DATA_55_const_net_31;
wire   [7:0]     TX_DATA_56_const_net_31;
wire   [7:0]     TX_DATA_57_const_net_31;
wire   [7:0]     TX_DATA_58_const_net_31;
wire   [7:0]     TX_DATA_59_const_net_31;
wire   [7:0]     TX_DATA_60_const_net_31;
wire   [7:0]     TX_DATA_61_const_net_31;
wire   [7:0]     TX_DATA_62_const_net_31;
wire   [7:0]     TX_DATA_63_const_net_31;
wire   [7:0]     TX_DATA_64_const_net_31;
wire   [7:0]     TX_DATA_65_const_net_31;
wire   [7:0]     TX_DATA_66_const_net_31;
wire   [7:0]     TX_DATA_67_const_net_31;
wire   [7:0]     TX_DATA_68_const_net_31;
wire   [7:0]     TX_DATA_69_const_net_31;
wire   [7:0]     TX_DATA_70_const_net_31;
wire   [7:0]     TX_DATA_71_const_net_31;
wire   [7:0]     TX_DATA_72_const_net_31;
wire   [7:0]     TX_DATA_73_const_net_31;
wire   [7:0]     TX_DATA_74_const_net_31;
wire   [7:0]     TX_DATA_75_const_net_31;
wire   [7:0]     TX_DATA_76_const_net_31;
wire   [7:0]     TX_DATA_77_const_net_31;
wire   [7:0]     TX_DATA_78_const_net_31;
wire   [7:0]     TX_DATA_79_const_net_31;
wire   [7:0]     TX_DATA_80_const_net_31;
wire   [7:0]     TX_DATA_81_const_net_31;
wire   [7:0]     TX_DATA_82_const_net_31;
wire   [7:0]     TX_DATA_83_const_net_31;
wire   [7:0]     TX_DATA_84_const_net_31;
wire   [7:0]     TX_DATA_85_const_net_31;
wire   [7:0]     TX_DATA_86_const_net_31;
wire   [7:0]     TX_DATA_87_const_net_31;
wire   [7:0]     TX_DATA_88_const_net_31;
wire   [7:0]     TX_DATA_89_const_net_31;
wire   [7:0]     TX_DATA_90_const_net_31;
wire   [7:0]     TX_DATA_91_const_net_31;
wire   [7:0]     TX_DATA_92_const_net_31;
wire   [7:0]     TX_DATA_93_const_net_31;
wire   [7:0]     TX_DATA_94_const_net_31;
wire   [7:0]     TX_DATA_95_const_net_31;
wire   [7:0]     TX_DATA_96_const_net_31;
wire   [7:0]     TX_DATA_97_const_net_31;
wire   [7:0]     TX_DATA_98_const_net_31;
wire   [7:0]     TX_DATA_99_const_net_31;
wire   [7:0]     TX_DATA_100_const_net_31;
wire   [7:0]     TX_DATA_101_const_net_31;
wire   [7:0]     TX_DATA_102_const_net_31;
wire   [7:0]     TX_DATA_103_const_net_31;
wire   [7:0]     TX_DATA_104_const_net_31;
wire   [7:0]     TX_DATA_105_const_net_31;
wire   [7:0]     TX_DATA_106_const_net_31;
wire   [7:0]     TX_DATA_107_const_net_31;
wire   [7:0]     TX_DATA_108_const_net_31;
wire   [7:0]     TX_DATA_109_const_net_31;
wire   [7:0]     TX_DATA_110_const_net_31;
wire   [7:0]     TX_DATA_111_const_net_31;
wire   [7:0]     TX_DATA_112_const_net_31;
wire   [7:0]     TX_DATA_113_const_net_31;
wire   [7:0]     TX_DATA_114_const_net_31;
wire   [7:0]     TX_DATA_115_const_net_31;
wire   [7:0]     TX_DATA_116_const_net_31;
wire   [7:0]     TX_DATA_117_const_net_31;
wire   [7:0]     TX_DATA_118_const_net_31;
wire   [7:0]     TX_DATA_119_const_net_31;
wire   [7:0]     TX_DATA_120_const_net_31;
wire   [7:0]     TX_DATA_121_const_net_31;
wire   [7:0]     TX_DATA_122_const_net_31;
wire   [7:0]     TX_DATA_123_const_net_31;
wire   [7:0]     TX_DATA_124_const_net_31;
wire   [7:0]     TX_DATA_125_const_net_31;
wire   [7:0]     TX_DATA_126_const_net_31;
wire   [7:0]     TX_DATA_127_const_net_31;
wire   [3:0]     OE_DATA_8_const_net_31;
wire   [3:0]     OE_DATA_9_const_net_31;
wire   [3:0]     OE_DATA_10_const_net_31;
wire   [3:0]     OE_DATA_11_const_net_31;
wire   [3:0]     OE_DATA_12_const_net_31;
wire   [3:0]     OE_DATA_13_const_net_31;
wire   [3:0]     OE_DATA_14_const_net_31;
wire   [3:0]     OE_DATA_15_const_net_31;
wire   [3:0]     OE_DATA_16_const_net_31;
wire   [3:0]     OE_DATA_17_const_net_31;
wire   [3:0]     OE_DATA_18_const_net_31;
wire   [3:0]     OE_DATA_19_const_net_31;
wire   [3:0]     OE_DATA_20_const_net_31;
wire   [3:0]     OE_DATA_21_const_net_31;
wire   [3:0]     OE_DATA_22_const_net_31;
wire   [3:0]     OE_DATA_23_const_net_31;
wire   [3:0]     OE_DATA_24_const_net_31;
wire   [3:0]     OE_DATA_25_const_net_31;
wire   [3:0]     OE_DATA_26_const_net_31;
wire   [3:0]     OE_DATA_27_const_net_31;
wire   [3:0]     OE_DATA_28_const_net_31;
wire   [3:0]     OE_DATA_29_const_net_31;
wire   [3:0]     OE_DATA_30_const_net_31;
wire   [3:0]     OE_DATA_31_const_net_31;
wire   [3:0]     OE_DATA_32_const_net_31;
wire   [3:0]     OE_DATA_33_const_net_31;
wire   [3:0]     OE_DATA_34_const_net_31;
wire   [3:0]     OE_DATA_35_const_net_31;
wire   [3:0]     OE_DATA_36_const_net_31;
wire   [3:0]     OE_DATA_37_const_net_31;
wire   [3:0]     OE_DATA_38_const_net_31;
wire   [3:0]     OE_DATA_39_const_net_31;
wire   [3:0]     OE_DATA_40_const_net_31;
wire   [3:0]     OE_DATA_41_const_net_31;
wire   [3:0]     OE_DATA_42_const_net_31;
wire   [3:0]     OE_DATA_43_const_net_31;
wire   [3:0]     OE_DATA_44_const_net_31;
wire   [3:0]     OE_DATA_45_const_net_31;
wire   [3:0]     OE_DATA_46_const_net_31;
wire   [3:0]     OE_DATA_47_const_net_31;
wire   [3:0]     OE_DATA_48_const_net_31;
wire   [3:0]     OE_DATA_49_const_net_31;
wire   [3:0]     OE_DATA_50_const_net_31;
wire   [3:0]     OE_DATA_51_const_net_31;
wire   [3:0]     OE_DATA_52_const_net_31;
wire   [3:0]     OE_DATA_53_const_net_31;
wire   [3:0]     OE_DATA_54_const_net_31;
wire   [3:0]     OE_DATA_55_const_net_31;
wire   [3:0]     OE_DATA_56_const_net_31;
wire   [3:0]     OE_DATA_57_const_net_31;
wire   [3:0]     OE_DATA_58_const_net_31;
wire   [3:0]     OE_DATA_59_const_net_31;
wire   [3:0]     OE_DATA_60_const_net_31;
wire   [3:0]     OE_DATA_61_const_net_31;
wire   [3:0]     OE_DATA_62_const_net_31;
wire   [3:0]     OE_DATA_63_const_net_31;
wire   [3:0]     OE_DATA_64_const_net_31;
wire   [3:0]     OE_DATA_65_const_net_31;
wire   [3:0]     OE_DATA_66_const_net_31;
wire   [3:0]     OE_DATA_67_const_net_31;
wire   [3:0]     OE_DATA_68_const_net_31;
wire   [3:0]     OE_DATA_69_const_net_31;
wire   [3:0]     OE_DATA_70_const_net_31;
wire   [3:0]     OE_DATA_71_const_net_31;
wire   [3:0]     OE_DATA_72_const_net_31;
wire   [3:0]     OE_DATA_73_const_net_31;
wire   [3:0]     OE_DATA_74_const_net_31;
wire   [3:0]     OE_DATA_75_const_net_31;
wire   [3:0]     OE_DATA_76_const_net_31;
wire   [3:0]     OE_DATA_77_const_net_31;
wire   [3:0]     OE_DATA_78_const_net_31;
wire   [3:0]     OE_DATA_79_const_net_31;
wire   [3:0]     OE_DATA_80_const_net_31;
wire   [3:0]     OE_DATA_81_const_net_31;
wire   [3:0]     OE_DATA_82_const_net_31;
wire   [3:0]     OE_DATA_83_const_net_31;
wire   [3:0]     OE_DATA_84_const_net_31;
wire   [3:0]     OE_DATA_85_const_net_31;
wire   [3:0]     OE_DATA_86_const_net_31;
wire   [3:0]     OE_DATA_87_const_net_31;
wire   [3:0]     OE_DATA_88_const_net_31;
wire   [3:0]     OE_DATA_89_const_net_31;
wire   [3:0]     OE_DATA_90_const_net_31;
wire   [3:0]     OE_DATA_91_const_net_31;
wire   [3:0]     OE_DATA_92_const_net_31;
wire   [3:0]     OE_DATA_93_const_net_31;
wire   [3:0]     OE_DATA_94_const_net_31;
wire   [3:0]     OE_DATA_95_const_net_31;
wire   [3:0]     OE_DATA_96_const_net_31;
wire   [3:0]     OE_DATA_97_const_net_31;
wire   [3:0]     OE_DATA_98_const_net_31;
wire   [3:0]     OE_DATA_99_const_net_31;
wire   [3:0]     OE_DATA_100_const_net_31;
wire   [3:0]     OE_DATA_101_const_net_31;
wire   [3:0]     OE_DATA_102_const_net_31;
wire   [3:0]     OE_DATA_103_const_net_31;
wire   [3:0]     OE_DATA_104_const_net_31;
wire   [3:0]     OE_DATA_105_const_net_31;
wire   [3:0]     OE_DATA_106_const_net_31;
wire   [3:0]     OE_DATA_107_const_net_31;
wire   [3:0]     OE_DATA_108_const_net_31;
wire   [3:0]     OE_DATA_109_const_net_31;
wire   [3:0]     OE_DATA_110_const_net_31;
wire   [3:0]     OE_DATA_111_const_net_31;
wire   [3:0]     OE_DATA_112_const_net_31;
wire   [3:0]     OE_DATA_113_const_net_31;
wire   [3:0]     OE_DATA_114_const_net_31;
wire   [3:0]     OE_DATA_115_const_net_31;
wire   [3:0]     OE_DATA_116_const_net_31;
wire   [3:0]     OE_DATA_117_const_net_31;
wire   [3:0]     OE_DATA_118_const_net_31;
wire   [3:0]     OE_DATA_119_const_net_31;
wire   [3:0]     OE_DATA_120_const_net_31;
wire   [3:0]     OE_DATA_121_const_net_31;
wire   [3:0]     OE_DATA_122_const_net_31;
wire   [3:0]     OE_DATA_123_const_net_31;
wire   [3:0]     OE_DATA_124_const_net_31;
wire   [3:0]     OE_DATA_125_const_net_31;
wire   [3:0]     OE_DATA_126_const_net_31;
wire   [3:0]     OE_DATA_127_const_net_31;
wire   [7:0]     PAD_I_const_net_6;
wire   [7:0]     PAD_N_const_net_6;
wire   [7:0]     PAD_I_N_const_net_6;
wire   [7:0]     TX_DATA_1_const_net_25;
wire   [7:0]     TX_DATA_2_const_net_27;
wire   [7:0]     TX_DATA_3_const_net_27;
wire   [7:0]     TX_DATA_4_const_net_27;
wire   [7:0]     TX_DATA_5_const_net_27;
wire   [7:0]     TX_DATA_6_const_net_27;
wire   [7:0]     TX_DATA_7_const_net_27;
wire   [7:0]     TX_DATA_8_const_net_31;
wire   [7:0]     TX_DATA_9_const_net_31;
wire   [7:0]     TX_DATA_10_const_net_31;
wire   [7:0]     TX_DATA_11_const_net_31;
wire   [7:0]     TX_DATA_12_const_net_32;
wire   [7:0]     TX_DATA_13_const_net_32;
wire   [7:0]     TX_DATA_14_const_net_32;
wire   [7:0]     TX_DATA_15_const_net_32;
wire   [7:0]     TX_DATA_16_const_net_32;
wire   [7:0]     TX_DATA_17_const_net_32;
wire   [7:0]     TX_DATA_18_const_net_32;
wire   [7:0]     TX_DATA_19_const_net_32;
wire   [7:0]     TX_DATA_20_const_net_32;
wire   [7:0]     TX_DATA_21_const_net_32;
wire   [7:0]     TX_DATA_22_const_net_32;
wire   [7:0]     TX_DATA_23_const_net_32;
wire   [7:0]     TX_DATA_24_const_net_32;
wire   [7:0]     TX_DATA_25_const_net_32;
wire   [7:0]     TX_DATA_26_const_net_32;
wire   [7:0]     TX_DATA_27_const_net_32;
wire   [7:0]     TX_DATA_28_const_net_32;
wire   [7:0]     TX_DATA_29_const_net_32;
wire   [7:0]     TX_DATA_30_const_net_32;
wire   [7:0]     TX_DATA_31_const_net_32;
wire   [7:0]     TX_DATA_32_const_net_32;
wire   [7:0]     TX_DATA_33_const_net_32;
wire   [7:0]     TX_DATA_34_const_net_32;
wire   [7:0]     TX_DATA_35_const_net_32;
wire   [7:0]     TX_DATA_36_const_net_32;
wire   [7:0]     TX_DATA_37_const_net_32;
wire   [7:0]     TX_DATA_38_const_net_32;
wire   [7:0]     TX_DATA_39_const_net_32;
wire   [7:0]     TX_DATA_40_const_net_32;
wire   [7:0]     TX_DATA_41_const_net_32;
wire   [7:0]     TX_DATA_42_const_net_32;
wire   [7:0]     TX_DATA_43_const_net_32;
wire   [7:0]     TX_DATA_44_const_net_32;
wire   [7:0]     TX_DATA_45_const_net_32;
wire   [7:0]     TX_DATA_46_const_net_32;
wire   [7:0]     TX_DATA_47_const_net_32;
wire   [7:0]     TX_DATA_48_const_net_32;
wire   [7:0]     TX_DATA_49_const_net_32;
wire   [7:0]     TX_DATA_50_const_net_32;
wire   [7:0]     TX_DATA_51_const_net_32;
wire   [7:0]     TX_DATA_52_const_net_32;
wire   [7:0]     TX_DATA_53_const_net_32;
wire   [7:0]     TX_DATA_54_const_net_32;
wire   [7:0]     TX_DATA_55_const_net_32;
wire   [7:0]     TX_DATA_56_const_net_32;
wire   [7:0]     TX_DATA_57_const_net_32;
wire   [7:0]     TX_DATA_58_const_net_32;
wire   [7:0]     TX_DATA_59_const_net_32;
wire   [7:0]     TX_DATA_60_const_net_32;
wire   [7:0]     TX_DATA_61_const_net_32;
wire   [7:0]     TX_DATA_62_const_net_32;
wire   [7:0]     TX_DATA_63_const_net_32;
wire   [7:0]     TX_DATA_64_const_net_32;
wire   [7:0]     TX_DATA_65_const_net_32;
wire   [7:0]     TX_DATA_66_const_net_32;
wire   [7:0]     TX_DATA_67_const_net_32;
wire   [7:0]     TX_DATA_68_const_net_32;
wire   [7:0]     TX_DATA_69_const_net_32;
wire   [7:0]     TX_DATA_70_const_net_32;
wire   [7:0]     TX_DATA_71_const_net_32;
wire   [7:0]     TX_DATA_72_const_net_32;
wire   [7:0]     TX_DATA_73_const_net_32;
wire   [7:0]     TX_DATA_74_const_net_32;
wire   [7:0]     TX_DATA_75_const_net_32;
wire   [7:0]     TX_DATA_76_const_net_32;
wire   [7:0]     TX_DATA_77_const_net_32;
wire   [7:0]     TX_DATA_78_const_net_32;
wire   [7:0]     TX_DATA_79_const_net_32;
wire   [7:0]     TX_DATA_80_const_net_32;
wire   [7:0]     TX_DATA_81_const_net_32;
wire   [7:0]     TX_DATA_82_const_net_32;
wire   [7:0]     TX_DATA_83_const_net_32;
wire   [7:0]     TX_DATA_84_const_net_32;
wire   [7:0]     TX_DATA_85_const_net_32;
wire   [7:0]     TX_DATA_86_const_net_32;
wire   [7:0]     TX_DATA_87_const_net_32;
wire   [7:0]     TX_DATA_88_const_net_32;
wire   [7:0]     TX_DATA_89_const_net_32;
wire   [7:0]     TX_DATA_90_const_net_32;
wire   [7:0]     TX_DATA_91_const_net_32;
wire   [7:0]     TX_DATA_92_const_net_32;
wire   [7:0]     TX_DATA_93_const_net_32;
wire   [7:0]     TX_DATA_94_const_net_32;
wire   [7:0]     TX_DATA_95_const_net_32;
wire   [7:0]     TX_DATA_96_const_net_32;
wire   [7:0]     TX_DATA_97_const_net_32;
wire   [7:0]     TX_DATA_98_const_net_32;
wire   [7:0]     TX_DATA_99_const_net_32;
wire   [7:0]     TX_DATA_100_const_net_32;
wire   [7:0]     TX_DATA_101_const_net_32;
wire   [7:0]     TX_DATA_102_const_net_32;
wire   [7:0]     TX_DATA_103_const_net_32;
wire   [7:0]     TX_DATA_104_const_net_32;
wire   [7:0]     TX_DATA_105_const_net_32;
wire   [7:0]     TX_DATA_106_const_net_32;
wire   [7:0]     TX_DATA_107_const_net_32;
wire   [7:0]     TX_DATA_108_const_net_32;
wire   [7:0]     TX_DATA_109_const_net_32;
wire   [7:0]     TX_DATA_110_const_net_32;
wire   [7:0]     TX_DATA_111_const_net_32;
wire   [7:0]     TX_DATA_112_const_net_32;
wire   [7:0]     TX_DATA_113_const_net_32;
wire   [7:0]     TX_DATA_114_const_net_32;
wire   [7:0]     TX_DATA_115_const_net_32;
wire   [7:0]     TX_DATA_116_const_net_32;
wire   [7:0]     TX_DATA_117_const_net_32;
wire   [7:0]     TX_DATA_118_const_net_32;
wire   [7:0]     TX_DATA_119_const_net_32;
wire   [7:0]     TX_DATA_120_const_net_32;
wire   [7:0]     TX_DATA_121_const_net_32;
wire   [7:0]     TX_DATA_122_const_net_32;
wire   [7:0]     TX_DATA_123_const_net_32;
wire   [7:0]     TX_DATA_124_const_net_32;
wire   [7:0]     TX_DATA_125_const_net_32;
wire   [7:0]     TX_DATA_126_const_net_32;
wire   [7:0]     TX_DATA_127_const_net_32;
wire   [3:0]     OE_DATA_1_const_net_28;
wire   [3:0]     OE_DATA_2_const_net_28;
wire   [3:0]     OE_DATA_3_const_net_28;
wire   [3:0]     OE_DATA_4_const_net_28;
wire   [3:0]     OE_DATA_5_const_net_28;
wire   [3:0]     OE_DATA_6_const_net_28;
wire   [3:0]     OE_DATA_7_const_net_28;
wire   [3:0]     OE_DATA_8_const_net_32;
wire   [3:0]     OE_DATA_9_const_net_32;
wire   [3:0]     OE_DATA_10_const_net_32;
wire   [3:0]     OE_DATA_11_const_net_32;
wire   [3:0]     OE_DATA_12_const_net_32;
wire   [3:0]     OE_DATA_13_const_net_32;
wire   [3:0]     OE_DATA_14_const_net_32;
wire   [3:0]     OE_DATA_15_const_net_32;
wire   [3:0]     OE_DATA_16_const_net_32;
wire   [3:0]     OE_DATA_17_const_net_32;
wire   [3:0]     OE_DATA_18_const_net_32;
wire   [3:0]     OE_DATA_19_const_net_32;
wire   [3:0]     OE_DATA_20_const_net_32;
wire   [3:0]     OE_DATA_21_const_net_32;
wire   [3:0]     OE_DATA_22_const_net_32;
wire   [3:0]     OE_DATA_23_const_net_32;
wire   [3:0]     OE_DATA_24_const_net_32;
wire   [3:0]     OE_DATA_25_const_net_32;
wire   [3:0]     OE_DATA_26_const_net_32;
wire   [3:0]     OE_DATA_27_const_net_32;
wire   [3:0]     OE_DATA_28_const_net_32;
wire   [3:0]     OE_DATA_29_const_net_32;
wire   [3:0]     OE_DATA_30_const_net_32;
wire   [3:0]     OE_DATA_31_const_net_32;
wire   [3:0]     OE_DATA_32_const_net_32;
wire   [3:0]     OE_DATA_33_const_net_32;
wire   [3:0]     OE_DATA_34_const_net_32;
wire   [3:0]     OE_DATA_35_const_net_32;
wire   [3:0]     OE_DATA_36_const_net_32;
wire   [3:0]     OE_DATA_37_const_net_32;
wire   [3:0]     OE_DATA_38_const_net_32;
wire   [3:0]     OE_DATA_39_const_net_32;
wire   [3:0]     OE_DATA_40_const_net_32;
wire   [3:0]     OE_DATA_41_const_net_32;
wire   [3:0]     OE_DATA_42_const_net_32;
wire   [3:0]     OE_DATA_43_const_net_32;
wire   [3:0]     OE_DATA_44_const_net_32;
wire   [3:0]     OE_DATA_45_const_net_32;
wire   [3:0]     OE_DATA_46_const_net_32;
wire   [3:0]     OE_DATA_47_const_net_32;
wire   [3:0]     OE_DATA_48_const_net_32;
wire   [3:0]     OE_DATA_49_const_net_32;
wire   [3:0]     OE_DATA_50_const_net_32;
wire   [3:0]     OE_DATA_51_const_net_32;
wire   [3:0]     OE_DATA_52_const_net_32;
wire   [3:0]     OE_DATA_53_const_net_32;
wire   [3:0]     OE_DATA_54_const_net_32;
wire   [3:0]     OE_DATA_55_const_net_32;
wire   [3:0]     OE_DATA_56_const_net_32;
wire   [3:0]     OE_DATA_57_const_net_32;
wire   [3:0]     OE_DATA_58_const_net_32;
wire   [3:0]     OE_DATA_59_const_net_32;
wire   [3:0]     OE_DATA_60_const_net_32;
wire   [3:0]     OE_DATA_61_const_net_32;
wire   [3:0]     OE_DATA_62_const_net_32;
wire   [3:0]     OE_DATA_63_const_net_32;
wire   [3:0]     OE_DATA_64_const_net_32;
wire   [3:0]     OE_DATA_65_const_net_32;
wire   [3:0]     OE_DATA_66_const_net_32;
wire   [3:0]     OE_DATA_67_const_net_32;
wire   [3:0]     OE_DATA_68_const_net_32;
wire   [3:0]     OE_DATA_69_const_net_32;
wire   [3:0]     OE_DATA_70_const_net_32;
wire   [3:0]     OE_DATA_71_const_net_32;
wire   [3:0]     OE_DATA_72_const_net_32;
wire   [3:0]     OE_DATA_73_const_net_32;
wire   [3:0]     OE_DATA_74_const_net_32;
wire   [3:0]     OE_DATA_75_const_net_32;
wire   [3:0]     OE_DATA_76_const_net_32;
wire   [3:0]     OE_DATA_77_const_net_32;
wire   [3:0]     OE_DATA_78_const_net_32;
wire   [3:0]     OE_DATA_79_const_net_32;
wire   [3:0]     OE_DATA_80_const_net_32;
wire   [3:0]     OE_DATA_81_const_net_32;
wire   [3:0]     OE_DATA_82_const_net_32;
wire   [3:0]     OE_DATA_83_const_net_32;
wire   [3:0]     OE_DATA_84_const_net_32;
wire   [3:0]     OE_DATA_85_const_net_32;
wire   [3:0]     OE_DATA_86_const_net_32;
wire   [3:0]     OE_DATA_87_const_net_32;
wire   [3:0]     OE_DATA_88_const_net_32;
wire   [3:0]     OE_DATA_89_const_net_32;
wire   [3:0]     OE_DATA_90_const_net_32;
wire   [3:0]     OE_DATA_91_const_net_32;
wire   [3:0]     OE_DATA_92_const_net_32;
wire   [3:0]     OE_DATA_93_const_net_32;
wire   [3:0]     OE_DATA_94_const_net_32;
wire   [3:0]     OE_DATA_95_const_net_32;
wire   [3:0]     OE_DATA_96_const_net_32;
wire   [3:0]     OE_DATA_97_const_net_32;
wire   [3:0]     OE_DATA_98_const_net_32;
wire   [3:0]     OE_DATA_99_const_net_32;
wire   [3:0]     OE_DATA_100_const_net_32;
wire   [3:0]     OE_DATA_101_const_net_32;
wire   [3:0]     OE_DATA_102_const_net_32;
wire   [3:0]     OE_DATA_103_const_net_32;
wire   [3:0]     OE_DATA_104_const_net_32;
wire   [3:0]     OE_DATA_105_const_net_32;
wire   [3:0]     OE_DATA_106_const_net_32;
wire   [3:0]     OE_DATA_107_const_net_32;
wire   [3:0]     OE_DATA_108_const_net_32;
wire   [3:0]     OE_DATA_109_const_net_32;
wire   [3:0]     OE_DATA_110_const_net_32;
wire   [3:0]     OE_DATA_111_const_net_32;
wire   [3:0]     OE_DATA_112_const_net_32;
wire   [3:0]     OE_DATA_113_const_net_32;
wire   [3:0]     OE_DATA_114_const_net_32;
wire   [3:0]     OE_DATA_115_const_net_32;
wire   [3:0]     OE_DATA_116_const_net_32;
wire   [3:0]     OE_DATA_117_const_net_32;
wire   [3:0]     OE_DATA_118_const_net_32;
wire   [3:0]     OE_DATA_119_const_net_32;
wire   [3:0]     OE_DATA_120_const_net_32;
wire   [3:0]     OE_DATA_121_const_net_32;
wire   [3:0]     OE_DATA_122_const_net_32;
wire   [3:0]     OE_DATA_123_const_net_32;
wire   [3:0]     OE_DATA_124_const_net_32;
wire   [3:0]     OE_DATA_125_const_net_32;
wire   [3:0]     OE_DATA_126_const_net_32;
wire   [3:0]     OE_DATA_127_const_net_32;
wire   [1:0]     RX_DQS_90_const_net_21;
wire   [2:0]     FIFO_WR_PTR_const_net_22;
wire   [2:0]     FIFO_RD_PTR_const_net_22;
wire   [2:0]     EYE_MONITOR_LANE_WIDTH_const_net_25;
wire   [1:0]     TX_DATA_1_const_net_26;
wire   [1:0]     TX_DATA_2_const_net_28;
wire   [1:0]     TX_DATA_3_const_net_28;
wire   [1:0]     TX_DATA_4_const_net_28;
wire   [1:0]     TX_DATA_5_const_net_28;
wire   [1:0]     TX_DATA_6_const_net_28;
wire   [1:0]     TX_DATA_7_const_net_28;
wire   [1:0]     TX_DATA_8_const_net_32;
wire   [1:0]     TX_DATA_9_const_net_32;
wire   [1:0]     TX_DATA_10_const_net_32;
wire   [1:0]     TX_DATA_11_const_net_32;
wire   [1:0]     TX_DATA_12_const_net_33;
wire   [1:0]     TX_DATA_13_const_net_33;
wire   [1:0]     TX_DATA_14_const_net_33;
wire   [1:0]     TX_DATA_15_const_net_33;
wire   [1:0]     TX_DATA_16_const_net_33;
wire   [1:0]     TX_DATA_17_const_net_33;
wire   [1:0]     TX_DATA_18_const_net_33;
wire   [1:0]     TX_DATA_19_const_net_33;
wire   [1:0]     TX_DATA_20_const_net_33;
wire   [1:0]     TX_DATA_21_const_net_33;
wire   [1:0]     TX_DATA_22_const_net_33;
wire   [1:0]     TX_DATA_23_const_net_33;
wire   [1:0]     TX_DATA_24_const_net_33;
wire   [1:0]     TX_DATA_25_const_net_33;
wire   [1:0]     TX_DATA_26_const_net_33;
wire   [1:0]     TX_DATA_27_const_net_33;
wire   [1:0]     TX_DATA_28_const_net_33;
wire   [1:0]     TX_DATA_29_const_net_33;
wire   [1:0]     TX_DATA_30_const_net_33;
wire   [1:0]     TX_DATA_31_const_net_33;
wire   [1:0]     TX_DATA_32_const_net_33;
wire   [1:0]     TX_DATA_33_const_net_33;
wire   [1:0]     TX_DATA_34_const_net_33;
wire   [1:0]     TX_DATA_35_const_net_33;
wire   [1:0]     TX_DATA_36_const_net_33;
wire   [1:0]     TX_DATA_37_const_net_33;
wire   [1:0]     TX_DATA_38_const_net_33;
wire   [1:0]     TX_DATA_39_const_net_33;
wire   [1:0]     TX_DATA_40_const_net_33;
wire   [1:0]     TX_DATA_41_const_net_33;
wire   [1:0]     TX_DATA_42_const_net_33;
wire   [1:0]     TX_DATA_43_const_net_33;
wire   [1:0]     TX_DATA_44_const_net_33;
wire   [1:0]     TX_DATA_45_const_net_33;
wire   [1:0]     TX_DATA_46_const_net_33;
wire   [1:0]     TX_DATA_47_const_net_33;
wire   [1:0]     TX_DATA_48_const_net_33;
wire   [1:0]     TX_DATA_49_const_net_33;
wire   [1:0]     TX_DATA_50_const_net_33;
wire   [1:0]     TX_DATA_51_const_net_33;
wire   [1:0]     TX_DATA_52_const_net_33;
wire   [1:0]     TX_DATA_53_const_net_33;
wire   [1:0]     TX_DATA_54_const_net_33;
wire   [1:0]     TX_DATA_55_const_net_33;
wire   [1:0]     TX_DATA_56_const_net_33;
wire   [1:0]     TX_DATA_57_const_net_33;
wire   [1:0]     TX_DATA_58_const_net_33;
wire   [1:0]     TX_DATA_59_const_net_33;
wire   [1:0]     TX_DATA_60_const_net_33;
wire   [1:0]     TX_DATA_61_const_net_33;
wire   [1:0]     TX_DATA_62_const_net_33;
wire   [1:0]     TX_DATA_63_const_net_33;
wire   [1:0]     TX_DATA_64_const_net_33;
wire   [1:0]     TX_DATA_65_const_net_33;
wire   [1:0]     TX_DATA_66_const_net_33;
wire   [1:0]     TX_DATA_67_const_net_33;
wire   [1:0]     TX_DATA_68_const_net_33;
wire   [1:0]     TX_DATA_69_const_net_33;
wire   [1:0]     TX_DATA_70_const_net_33;
wire   [1:0]     TX_DATA_71_const_net_33;
wire   [1:0]     TX_DATA_72_const_net_33;
wire   [1:0]     TX_DATA_73_const_net_33;
wire   [1:0]     TX_DATA_74_const_net_33;
wire   [1:0]     TX_DATA_75_const_net_33;
wire   [1:0]     TX_DATA_76_const_net_33;
wire   [1:0]     TX_DATA_77_const_net_33;
wire   [1:0]     TX_DATA_78_const_net_33;
wire   [1:0]     TX_DATA_79_const_net_33;
wire   [1:0]     TX_DATA_80_const_net_33;
wire   [1:0]     TX_DATA_81_const_net_33;
wire   [1:0]     TX_DATA_82_const_net_33;
wire   [1:0]     TX_DATA_83_const_net_33;
wire   [1:0]     TX_DATA_84_const_net_33;
wire   [1:0]     TX_DATA_85_const_net_33;
wire   [1:0]     TX_DATA_86_const_net_33;
wire   [1:0]     TX_DATA_87_const_net_33;
wire   [1:0]     TX_DATA_88_const_net_33;
wire   [1:0]     TX_DATA_89_const_net_33;
wire   [1:0]     TX_DATA_90_const_net_33;
wire   [1:0]     TX_DATA_91_const_net_33;
wire   [1:0]     TX_DATA_92_const_net_33;
wire   [1:0]     TX_DATA_93_const_net_33;
wire   [1:0]     TX_DATA_94_const_net_33;
wire   [1:0]     TX_DATA_95_const_net_33;
wire   [1:0]     TX_DATA_96_const_net_33;
wire   [1:0]     TX_DATA_97_const_net_33;
wire   [1:0]     TX_DATA_98_const_net_33;
wire   [1:0]     TX_DATA_99_const_net_33;
wire   [1:0]     TX_DATA_100_const_net_33;
wire   [1:0]     TX_DATA_101_const_net_33;
wire   [1:0]     TX_DATA_102_const_net_33;
wire   [1:0]     TX_DATA_103_const_net_33;
wire   [1:0]     TX_DATA_104_const_net_33;
wire   [1:0]     TX_DATA_105_const_net_33;
wire   [1:0]     TX_DATA_106_const_net_33;
wire   [1:0]     TX_DATA_107_const_net_33;
wire   [1:0]     TX_DATA_108_const_net_33;
wire   [1:0]     TX_DATA_109_const_net_33;
wire   [1:0]     TX_DATA_110_const_net_33;
wire   [1:0]     TX_DATA_111_const_net_33;
wire   [1:0]     TX_DATA_112_const_net_33;
wire   [1:0]     TX_DATA_113_const_net_33;
wire   [1:0]     TX_DATA_114_const_net_33;
wire   [1:0]     TX_DATA_115_const_net_33;
wire   [1:0]     TX_DATA_116_const_net_33;
wire   [1:0]     TX_DATA_117_const_net_33;
wire   [1:0]     TX_DATA_118_const_net_33;
wire   [1:0]     TX_DATA_119_const_net_33;
wire   [1:0]     TX_DATA_120_const_net_33;
wire   [1:0]     TX_DATA_121_const_net_33;
wire   [1:0]     TX_DATA_122_const_net_33;
wire   [1:0]     TX_DATA_123_const_net_33;
wire   [1:0]     TX_DATA_124_const_net_33;
wire   [1:0]     TX_DATA_125_const_net_33;
wire   [1:0]     TX_DATA_126_const_net_33;
wire   [1:0]     TX_DATA_127_const_net_33;
wire   [1:0]     OE_DATA_1_const_net_29;
wire   [1:0]     OE_DATA_2_const_net_29;
wire   [1:0]     OE_DATA_3_const_net_29;
wire   [1:0]     OE_DATA_4_const_net_29;
wire   [1:0]     OE_DATA_5_const_net_29;
wire   [1:0]     OE_DATA_6_const_net_29;
wire   [1:0]     OE_DATA_7_const_net_29;
wire   [1:0]     OE_DATA_8_const_net_33;
wire   [1:0]     OE_DATA_9_const_net_33;
wire   [1:0]     OE_DATA_10_const_net_33;
wire   [1:0]     OE_DATA_11_const_net_33;
wire   [1:0]     OE_DATA_12_const_net_33;
wire   [1:0]     OE_DATA_13_const_net_33;
wire   [1:0]     OE_DATA_14_const_net_33;
wire   [1:0]     OE_DATA_15_const_net_33;
wire   [1:0]     OE_DATA_16_const_net_33;
wire   [1:0]     OE_DATA_17_const_net_33;
wire   [1:0]     OE_DATA_18_const_net_33;
wire   [1:0]     OE_DATA_19_const_net_33;
wire   [1:0]     OE_DATA_20_const_net_33;
wire   [1:0]     OE_DATA_21_const_net_33;
wire   [1:0]     OE_DATA_22_const_net_33;
wire   [1:0]     OE_DATA_23_const_net_33;
wire   [1:0]     OE_DATA_24_const_net_33;
wire   [1:0]     OE_DATA_25_const_net_33;
wire   [1:0]     OE_DATA_26_const_net_33;
wire   [1:0]     OE_DATA_27_const_net_33;
wire   [1:0]     OE_DATA_28_const_net_33;
wire   [1:0]     OE_DATA_29_const_net_33;
wire   [1:0]     OE_DATA_30_const_net_33;
wire   [1:0]     OE_DATA_31_const_net_33;
wire   [1:0]     OE_DATA_32_const_net_33;
wire   [1:0]     OE_DATA_33_const_net_33;
wire   [1:0]     OE_DATA_34_const_net_33;
wire   [1:0]     OE_DATA_35_const_net_33;
wire   [1:0]     OE_DATA_36_const_net_33;
wire   [1:0]     OE_DATA_37_const_net_33;
wire   [1:0]     OE_DATA_38_const_net_33;
wire   [1:0]     OE_DATA_39_const_net_33;
wire   [1:0]     OE_DATA_40_const_net_33;
wire   [1:0]     OE_DATA_41_const_net_33;
wire   [1:0]     OE_DATA_42_const_net_33;
wire   [1:0]     OE_DATA_43_const_net_33;
wire   [1:0]     OE_DATA_44_const_net_33;
wire   [1:0]     OE_DATA_45_const_net_33;
wire   [1:0]     OE_DATA_46_const_net_33;
wire   [1:0]     OE_DATA_47_const_net_33;
wire   [1:0]     OE_DATA_48_const_net_33;
wire   [1:0]     OE_DATA_49_const_net_33;
wire   [1:0]     OE_DATA_50_const_net_33;
wire   [1:0]     OE_DATA_51_const_net_33;
wire   [1:0]     OE_DATA_52_const_net_33;
wire   [1:0]     OE_DATA_53_const_net_33;
wire   [1:0]     OE_DATA_54_const_net_33;
wire   [1:0]     OE_DATA_55_const_net_33;
wire   [1:0]     OE_DATA_56_const_net_33;
wire   [1:0]     OE_DATA_57_const_net_33;
wire   [1:0]     OE_DATA_58_const_net_33;
wire   [1:0]     OE_DATA_59_const_net_33;
wire   [1:0]     OE_DATA_60_const_net_33;
wire   [1:0]     OE_DATA_61_const_net_33;
wire   [1:0]     OE_DATA_62_const_net_33;
wire   [1:0]     OE_DATA_63_const_net_33;
wire   [1:0]     OE_DATA_64_const_net_33;
wire   [1:0]     OE_DATA_65_const_net_33;
wire   [1:0]     OE_DATA_66_const_net_33;
wire   [1:0]     OE_DATA_67_const_net_33;
wire   [1:0]     OE_DATA_68_const_net_33;
wire   [1:0]     OE_DATA_69_const_net_33;
wire   [1:0]     OE_DATA_70_const_net_33;
wire   [1:0]     OE_DATA_71_const_net_33;
wire   [1:0]     OE_DATA_72_const_net_33;
wire   [1:0]     OE_DATA_73_const_net_33;
wire   [1:0]     OE_DATA_74_const_net_33;
wire   [1:0]     OE_DATA_75_const_net_33;
wire   [1:0]     OE_DATA_76_const_net_33;
wire   [1:0]     OE_DATA_77_const_net_33;
wire   [1:0]     OE_DATA_78_const_net_33;
wire   [1:0]     OE_DATA_79_const_net_33;
wire   [1:0]     OE_DATA_80_const_net_33;
wire   [1:0]     OE_DATA_81_const_net_33;
wire   [1:0]     OE_DATA_82_const_net_33;
wire   [1:0]     OE_DATA_83_const_net_33;
wire   [1:0]     OE_DATA_84_const_net_33;
wire   [1:0]     OE_DATA_85_const_net_33;
wire   [1:0]     OE_DATA_86_const_net_33;
wire   [1:0]     OE_DATA_87_const_net_33;
wire   [1:0]     OE_DATA_88_const_net_33;
wire   [1:0]     OE_DATA_89_const_net_33;
wire   [1:0]     OE_DATA_90_const_net_33;
wire   [1:0]     OE_DATA_91_const_net_33;
wire   [1:0]     OE_DATA_92_const_net_33;
wire   [1:0]     OE_DATA_93_const_net_33;
wire   [1:0]     OE_DATA_94_const_net_33;
wire   [1:0]     OE_DATA_95_const_net_33;
wire   [1:0]     OE_DATA_96_const_net_33;
wire   [1:0]     OE_DATA_97_const_net_33;
wire   [1:0]     OE_DATA_98_const_net_33;
wire   [1:0]     OE_DATA_99_const_net_33;
wire   [1:0]     OE_DATA_100_const_net_33;
wire   [1:0]     OE_DATA_101_const_net_33;
wire   [1:0]     OE_DATA_102_const_net_33;
wire   [1:0]     OE_DATA_103_const_net_33;
wire   [1:0]     OE_DATA_104_const_net_33;
wire   [1:0]     OE_DATA_105_const_net_33;
wire   [1:0]     OE_DATA_106_const_net_33;
wire   [1:0]     OE_DATA_107_const_net_33;
wire   [1:0]     OE_DATA_108_const_net_33;
wire   [1:0]     OE_DATA_109_const_net_33;
wire   [1:0]     OE_DATA_110_const_net_33;
wire   [1:0]     OE_DATA_111_const_net_33;
wire   [1:0]     OE_DATA_112_const_net_33;
wire   [1:0]     OE_DATA_113_const_net_33;
wire   [1:0]     OE_DATA_114_const_net_33;
wire   [1:0]     OE_DATA_115_const_net_33;
wire   [1:0]     OE_DATA_116_const_net_33;
wire   [1:0]     OE_DATA_117_const_net_33;
wire   [1:0]     OE_DATA_118_const_net_33;
wire   [1:0]     OE_DATA_119_const_net_33;
wire   [1:0]     OE_DATA_120_const_net_33;
wire   [1:0]     OE_DATA_121_const_net_33;
wire   [1:0]     OE_DATA_122_const_net_33;
wire   [1:0]     OE_DATA_123_const_net_33;
wire   [1:0]     OE_DATA_124_const_net_33;
wire   [1:0]     OE_DATA_125_const_net_33;
wire   [1:0]     OE_DATA_126_const_net_33;
wire   [1:0]     OE_DATA_127_const_net_33;
wire   [1:0]     RX_DQS_90_const_net_22;
wire   [2:0]     EYE_MONITOR_LANE_WIDTH_const_net_26;
wire   [7:0]     TX_DATA_1_const_net_27;
wire   [7:0]     TX_DATA_2_const_net_29;
wire   [7:0]     TX_DATA_3_const_net_29;
wire   [7:0]     TX_DATA_4_const_net_29;
wire   [7:0]     TX_DATA_5_const_net_29;
wire   [7:0]     TX_DATA_6_const_net_29;
wire   [7:0]     TX_DATA_7_const_net_29;
wire   [7:0]     TX_DATA_8_const_net_33;
wire   [7:0]     TX_DATA_9_const_net_33;
wire   [7:0]     TX_DATA_10_const_net_33;
wire   [7:0]     TX_DATA_11_const_net_33;
wire   [7:0]     TX_DATA_12_const_net_34;
wire   [7:0]     TX_DATA_13_const_net_34;
wire   [7:0]     TX_DATA_14_const_net_34;
wire   [7:0]     TX_DATA_15_const_net_34;
wire   [7:0]     TX_DATA_16_const_net_34;
wire   [7:0]     TX_DATA_17_const_net_34;
wire   [7:0]     TX_DATA_18_const_net_34;
wire   [7:0]     TX_DATA_19_const_net_34;
wire   [7:0]     TX_DATA_20_const_net_34;
wire   [7:0]     TX_DATA_21_const_net_34;
wire   [7:0]     TX_DATA_22_const_net_34;
wire   [7:0]     TX_DATA_23_const_net_34;
wire   [7:0]     TX_DATA_24_const_net_34;
wire   [7:0]     TX_DATA_25_const_net_34;
wire   [7:0]     TX_DATA_26_const_net_34;
wire   [7:0]     TX_DATA_27_const_net_34;
wire   [7:0]     TX_DATA_28_const_net_34;
wire   [7:0]     TX_DATA_29_const_net_34;
wire   [7:0]     TX_DATA_30_const_net_34;
wire   [7:0]     TX_DATA_31_const_net_34;
wire   [7:0]     TX_DATA_32_const_net_34;
wire   [7:0]     TX_DATA_33_const_net_34;
wire   [7:0]     TX_DATA_34_const_net_34;
wire   [7:0]     TX_DATA_35_const_net_34;
wire   [7:0]     TX_DATA_36_const_net_34;
wire   [7:0]     TX_DATA_37_const_net_34;
wire   [7:0]     TX_DATA_38_const_net_34;
wire   [7:0]     TX_DATA_39_const_net_34;
wire   [7:0]     TX_DATA_40_const_net_34;
wire   [7:0]     TX_DATA_41_const_net_34;
wire   [7:0]     TX_DATA_42_const_net_34;
wire   [7:0]     TX_DATA_43_const_net_34;
wire   [7:0]     TX_DATA_44_const_net_34;
wire   [7:0]     TX_DATA_45_const_net_34;
wire   [7:0]     TX_DATA_46_const_net_34;
wire   [7:0]     TX_DATA_47_const_net_34;
wire   [7:0]     TX_DATA_48_const_net_34;
wire   [7:0]     TX_DATA_49_const_net_34;
wire   [7:0]     TX_DATA_50_const_net_34;
wire   [7:0]     TX_DATA_51_const_net_34;
wire   [7:0]     TX_DATA_52_const_net_34;
wire   [7:0]     TX_DATA_53_const_net_34;
wire   [7:0]     TX_DATA_54_const_net_34;
wire   [7:0]     TX_DATA_55_const_net_34;
wire   [7:0]     TX_DATA_56_const_net_34;
wire   [7:0]     TX_DATA_57_const_net_34;
wire   [7:0]     TX_DATA_58_const_net_34;
wire   [7:0]     TX_DATA_59_const_net_34;
wire   [7:0]     TX_DATA_60_const_net_34;
wire   [7:0]     TX_DATA_61_const_net_34;
wire   [7:0]     TX_DATA_62_const_net_34;
wire   [7:0]     TX_DATA_63_const_net_34;
wire   [7:0]     TX_DATA_64_const_net_34;
wire   [7:0]     TX_DATA_65_const_net_34;
wire   [7:0]     TX_DATA_66_const_net_34;
wire   [7:0]     TX_DATA_67_const_net_34;
wire   [7:0]     TX_DATA_68_const_net_34;
wire   [7:0]     TX_DATA_69_const_net_34;
wire   [7:0]     TX_DATA_70_const_net_34;
wire   [7:0]     TX_DATA_71_const_net_34;
wire   [7:0]     TX_DATA_72_const_net_34;
wire   [7:0]     TX_DATA_73_const_net_34;
wire   [7:0]     TX_DATA_74_const_net_34;
wire   [7:0]     TX_DATA_75_const_net_34;
wire   [7:0]     TX_DATA_76_const_net_34;
wire   [7:0]     TX_DATA_77_const_net_34;
wire   [7:0]     TX_DATA_78_const_net_34;
wire   [7:0]     TX_DATA_79_const_net_34;
wire   [7:0]     TX_DATA_80_const_net_34;
wire   [7:0]     TX_DATA_81_const_net_34;
wire   [7:0]     TX_DATA_82_const_net_34;
wire   [7:0]     TX_DATA_83_const_net_34;
wire   [7:0]     TX_DATA_84_const_net_34;
wire   [7:0]     TX_DATA_85_const_net_34;
wire   [7:0]     TX_DATA_86_const_net_34;
wire   [7:0]     TX_DATA_87_const_net_34;
wire   [7:0]     TX_DATA_88_const_net_34;
wire   [7:0]     TX_DATA_89_const_net_34;
wire   [7:0]     TX_DATA_90_const_net_34;
wire   [7:0]     TX_DATA_91_const_net_34;
wire   [7:0]     TX_DATA_92_const_net_34;
wire   [7:0]     TX_DATA_93_const_net_34;
wire   [7:0]     TX_DATA_94_const_net_34;
wire   [7:0]     TX_DATA_95_const_net_34;
wire   [7:0]     TX_DATA_96_const_net_34;
wire   [7:0]     TX_DATA_97_const_net_34;
wire   [7:0]     TX_DATA_98_const_net_34;
wire   [7:0]     TX_DATA_99_const_net_34;
wire   [7:0]     TX_DATA_100_const_net_34;
wire   [7:0]     TX_DATA_101_const_net_34;
wire   [7:0]     TX_DATA_102_const_net_34;
wire   [7:0]     TX_DATA_103_const_net_34;
wire   [7:0]     TX_DATA_104_const_net_34;
wire   [7:0]     TX_DATA_105_const_net_34;
wire   [7:0]     TX_DATA_106_const_net_34;
wire   [7:0]     TX_DATA_107_const_net_34;
wire   [7:0]     TX_DATA_108_const_net_34;
wire   [7:0]     TX_DATA_109_const_net_34;
wire   [7:0]     TX_DATA_110_const_net_34;
wire   [7:0]     TX_DATA_111_const_net_34;
wire   [7:0]     TX_DATA_112_const_net_34;
wire   [7:0]     TX_DATA_113_const_net_34;
wire   [7:0]     TX_DATA_114_const_net_34;
wire   [7:0]     TX_DATA_115_const_net_34;
wire   [7:0]     TX_DATA_116_const_net_34;
wire   [7:0]     TX_DATA_117_const_net_34;
wire   [7:0]     TX_DATA_118_const_net_34;
wire   [7:0]     TX_DATA_119_const_net_34;
wire   [7:0]     TX_DATA_120_const_net_34;
wire   [7:0]     TX_DATA_121_const_net_34;
wire   [7:0]     TX_DATA_122_const_net_34;
wire   [7:0]     TX_DATA_123_const_net_34;
wire   [7:0]     TX_DATA_124_const_net_34;
wire   [7:0]     TX_DATA_125_const_net_34;
wire   [7:0]     TX_DATA_126_const_net_34;
wire   [7:0]     TX_DATA_127_const_net_34;
wire   [3:0]     OE_DATA_1_const_net_30;
wire   [3:0]     OE_DATA_2_const_net_30;
wire   [3:0]     OE_DATA_3_const_net_30;
wire   [3:0]     OE_DATA_4_const_net_30;
wire   [3:0]     OE_DATA_5_const_net_30;
wire   [3:0]     OE_DATA_6_const_net_30;
wire   [3:0]     OE_DATA_7_const_net_30;
wire   [3:0]     OE_DATA_8_const_net_34;
wire   [3:0]     OE_DATA_9_const_net_34;
wire   [3:0]     OE_DATA_10_const_net_34;
wire   [3:0]     OE_DATA_11_const_net_34;
wire   [3:0]     OE_DATA_12_const_net_34;
wire   [3:0]     OE_DATA_13_const_net_34;
wire   [3:0]     OE_DATA_14_const_net_34;
wire   [3:0]     OE_DATA_15_const_net_34;
wire   [3:0]     OE_DATA_16_const_net_34;
wire   [3:0]     OE_DATA_17_const_net_34;
wire   [3:0]     OE_DATA_18_const_net_34;
wire   [3:0]     OE_DATA_19_const_net_34;
wire   [3:0]     OE_DATA_20_const_net_34;
wire   [3:0]     OE_DATA_21_const_net_34;
wire   [3:0]     OE_DATA_22_const_net_34;
wire   [3:0]     OE_DATA_23_const_net_34;
wire   [3:0]     OE_DATA_24_const_net_34;
wire   [3:0]     OE_DATA_25_const_net_34;
wire   [3:0]     OE_DATA_26_const_net_34;
wire   [3:0]     OE_DATA_27_const_net_34;
wire   [3:0]     OE_DATA_28_const_net_34;
wire   [3:0]     OE_DATA_29_const_net_34;
wire   [3:0]     OE_DATA_30_const_net_34;
wire   [3:0]     OE_DATA_31_const_net_34;
wire   [3:0]     OE_DATA_32_const_net_34;
wire   [3:0]     OE_DATA_33_const_net_34;
wire   [3:0]     OE_DATA_34_const_net_34;
wire   [3:0]     OE_DATA_35_const_net_34;
wire   [3:0]     OE_DATA_36_const_net_34;
wire   [3:0]     OE_DATA_37_const_net_34;
wire   [3:0]     OE_DATA_38_const_net_34;
wire   [3:0]     OE_DATA_39_const_net_34;
wire   [3:0]     OE_DATA_40_const_net_34;
wire   [3:0]     OE_DATA_41_const_net_34;
wire   [3:0]     OE_DATA_42_const_net_34;
wire   [3:0]     OE_DATA_43_const_net_34;
wire   [3:0]     OE_DATA_44_const_net_34;
wire   [3:0]     OE_DATA_45_const_net_34;
wire   [3:0]     OE_DATA_46_const_net_34;
wire   [3:0]     OE_DATA_47_const_net_34;
wire   [3:0]     OE_DATA_48_const_net_34;
wire   [3:0]     OE_DATA_49_const_net_34;
wire   [3:0]     OE_DATA_50_const_net_34;
wire   [3:0]     OE_DATA_51_const_net_34;
wire   [3:0]     OE_DATA_52_const_net_34;
wire   [3:0]     OE_DATA_53_const_net_34;
wire   [3:0]     OE_DATA_54_const_net_34;
wire   [3:0]     OE_DATA_55_const_net_34;
wire   [3:0]     OE_DATA_56_const_net_34;
wire   [3:0]     OE_DATA_57_const_net_34;
wire   [3:0]     OE_DATA_58_const_net_34;
wire   [3:0]     OE_DATA_59_const_net_34;
wire   [3:0]     OE_DATA_60_const_net_34;
wire   [3:0]     OE_DATA_61_const_net_34;
wire   [3:0]     OE_DATA_62_const_net_34;
wire   [3:0]     OE_DATA_63_const_net_34;
wire   [3:0]     OE_DATA_64_const_net_34;
wire   [3:0]     OE_DATA_65_const_net_34;
wire   [3:0]     OE_DATA_66_const_net_34;
wire   [3:0]     OE_DATA_67_const_net_34;
wire   [3:0]     OE_DATA_68_const_net_34;
wire   [3:0]     OE_DATA_69_const_net_34;
wire   [3:0]     OE_DATA_70_const_net_34;
wire   [3:0]     OE_DATA_71_const_net_34;
wire   [3:0]     OE_DATA_72_const_net_34;
wire   [3:0]     OE_DATA_73_const_net_34;
wire   [3:0]     OE_DATA_74_const_net_34;
wire   [3:0]     OE_DATA_75_const_net_34;
wire   [3:0]     OE_DATA_76_const_net_34;
wire   [3:0]     OE_DATA_77_const_net_34;
wire   [3:0]     OE_DATA_78_const_net_34;
wire   [3:0]     OE_DATA_79_const_net_34;
wire   [3:0]     OE_DATA_80_const_net_34;
wire   [3:0]     OE_DATA_81_const_net_34;
wire   [3:0]     OE_DATA_82_const_net_34;
wire   [3:0]     OE_DATA_83_const_net_34;
wire   [3:0]     OE_DATA_84_const_net_34;
wire   [3:0]     OE_DATA_85_const_net_34;
wire   [3:0]     OE_DATA_86_const_net_34;
wire   [3:0]     OE_DATA_87_const_net_34;
wire   [3:0]     OE_DATA_88_const_net_34;
wire   [3:0]     OE_DATA_89_const_net_34;
wire   [3:0]     OE_DATA_90_const_net_34;
wire   [3:0]     OE_DATA_91_const_net_34;
wire   [3:0]     OE_DATA_92_const_net_34;
wire   [3:0]     OE_DATA_93_const_net_34;
wire   [3:0]     OE_DATA_94_const_net_34;
wire   [3:0]     OE_DATA_95_const_net_34;
wire   [3:0]     OE_DATA_96_const_net_34;
wire   [3:0]     OE_DATA_97_const_net_34;
wire   [3:0]     OE_DATA_98_const_net_34;
wire   [3:0]     OE_DATA_99_const_net_34;
wire   [3:0]     OE_DATA_100_const_net_34;
wire   [3:0]     OE_DATA_101_const_net_34;
wire   [3:0]     OE_DATA_102_const_net_34;
wire   [3:0]     OE_DATA_103_const_net_34;
wire   [3:0]     OE_DATA_104_const_net_34;
wire   [3:0]     OE_DATA_105_const_net_34;
wire   [3:0]     OE_DATA_106_const_net_34;
wire   [3:0]     OE_DATA_107_const_net_34;
wire   [3:0]     OE_DATA_108_const_net_34;
wire   [3:0]     OE_DATA_109_const_net_34;
wire   [3:0]     OE_DATA_110_const_net_34;
wire   [3:0]     OE_DATA_111_const_net_34;
wire   [3:0]     OE_DATA_112_const_net_34;
wire   [3:0]     OE_DATA_113_const_net_34;
wire   [3:0]     OE_DATA_114_const_net_34;
wire   [3:0]     OE_DATA_115_const_net_34;
wire   [3:0]     OE_DATA_116_const_net_34;
wire   [3:0]     OE_DATA_117_const_net_34;
wire   [3:0]     OE_DATA_118_const_net_34;
wire   [3:0]     OE_DATA_119_const_net_34;
wire   [3:0]     OE_DATA_120_const_net_34;
wire   [3:0]     OE_DATA_121_const_net_34;
wire   [3:0]     OE_DATA_122_const_net_34;
wire   [3:0]     OE_DATA_123_const_net_34;
wire   [3:0]     OE_DATA_124_const_net_34;
wire   [3:0]     OE_DATA_125_const_net_34;
wire   [3:0]     OE_DATA_126_const_net_34;
wire   [3:0]     OE_DATA_127_const_net_34;
wire   [2:0]     READ_CLK_SEL_const_net_0;
wire   [2:0]     EYE_MONITOR_WIDTH_IN_const_net_4;
wire   [7:0]     CDR_CLK_A_SEL_const_net_0;
wire   [10:0]    CDR_CLK_B_SEL_const_net_4;
//--------------------------------------------------------------------
// Inverted Nets
//--------------------------------------------------------------------
wire             SYNC_SYS_RST_N_net_1;
wire             SYNC_SYS_RST_N_OUT_PRE_INV0_0;
//--------------------------------------------------------------------
// Constant assignments
//--------------------------------------------------------------------
assign DFI_CALVL_RESP_const_net_0          = 2'h0;
assign VCC_net                             = 1'b1;
assign GND_net                             = 1'b0;
assign DFI_PHYUPD_TYPE_const_net_0         = 2'h0;
assign OE_DATA_0_const_net_0               = 4'hF;
assign OE_DATA_1_const_net_0               = 4'hF;
assign OE_DATA_2_const_net_0               = 4'hF;
assign OE_DATA_3_const_net_0               = 4'hF;
assign OE_DATA_4_const_net_0               = 4'hF;
assign OE_DATA_5_const_net_0               = 4'hF;
assign OE_DATA_6_const_net_0               = 4'hF;
assign OE_DATA_7_const_net_0               = 4'hF;
assign OE_DATA_8_const_net_0               = 4'hF;
assign OE_DATA_9_const_net_0               = 4'hF;
assign OE_DATA_10_const_net_0              = 4'hF;
assign OE_DATA_11_const_net_0              = 4'hF;
assign OE_DATA_0_const_net_1               = 4'hF;
assign OE_DATA_0_const_net_2               = 4'hF;
assign OE_DATA_0_const_net_3               = 4'hF;
assign OE_DATA_1_const_net_1               = 4'hF;
assign OE_DATA_0_const_net_4               = 4'hF;
assign OE_DATA_1_const_net_2               = 4'hF;
assign OE_DATA_0_const_net_5               = 4'hF;
assign OE_DATA_0_const_net_6               = 4'hF;
assign OE_DATA_0_const_net_7               = 4'hF;
assign OE_DATA_0_const_net_8               = 4'hF;
assign OE_DATA_0_const_net_9               = 4'hF;
assign OE_DATA_0_const_net_10              = 4'hF;
assign TRAINING_PATTERN_const_net_0        = 8'hAA;
assign OE_DATA_0_const_net_11              = 4'hF;
assign EYE_MONITOR_WIDTH_IN_const_net_0    = 3'h2;
assign TX_DATA_0_const_net_0               = 8'h55;
assign TX_DATA_0_const_net_1               = 2'h0;
assign OE_DATA_0_const_net_12              = 2'h3;
assign EYE_MONITOR_WIDTH_IN_const_net_1    = 3'h2;
assign TX_DATA_0_const_net_2               = 8'h55;
assign TX_DATA_0_const_net_3               = 2'h0;
assign OE_DATA_0_const_net_13              = 2'h3;
assign EYE_MONITOR_WIDTH_IN_const_net_2    = 3'h2;
assign TX_DATA_0_const_net_4               = 8'h55;
assign TX_DATA_0_const_net_5               = 2'h0;
assign OE_DATA_0_const_net_14              = 2'h3;
assign EYE_MONITOR_WIDTH_IN_const_net_3    = 3'h2;
assign TX_DATA_0_const_net_6               = 8'h55;
assign TX_DATA_0_const_net_7               = 2'h0;
assign OE_DATA_0_const_net_15              = 2'h3;
assign RX_DQS_90_const_net_0               = 2'h0;
assign FIFO_WR_PTR_const_net_0             = 3'h0;
assign FIFO_RD_PTR_const_net_0             = 3'h0;
assign EYE_MONITOR_LANE_WIDTH_const_net_0  = 3'h0;
assign TX_DATA_12_const_net_0              = 4'h0;
assign TX_DATA_13_const_net_0              = 4'h0;
assign TX_DATA_14_const_net_0              = 4'h0;
assign TX_DATA_15_const_net_0              = 4'h0;
assign TX_DATA_16_const_net_0              = 4'h0;
assign TX_DATA_17_const_net_0              = 4'h0;
assign TX_DATA_18_const_net_0              = 4'h0;
assign TX_DATA_19_const_net_0              = 4'h0;
assign TX_DATA_20_const_net_0              = 4'h0;
assign TX_DATA_21_const_net_0              = 4'h0;
assign TX_DATA_22_const_net_0              = 4'h0;
assign TX_DATA_23_const_net_0              = 4'h0;
assign TX_DATA_24_const_net_0              = 4'h0;
assign TX_DATA_25_const_net_0              = 4'h0;
assign TX_DATA_26_const_net_0              = 4'h0;
assign TX_DATA_27_const_net_0              = 4'h0;
assign TX_DATA_28_const_net_0              = 4'h0;
assign TX_DATA_29_const_net_0              = 4'h0;
assign TX_DATA_30_const_net_0              = 4'h0;
assign TX_DATA_31_const_net_0              = 4'h0;
assign TX_DATA_32_const_net_0              = 4'h0;
assign TX_DATA_33_const_net_0              = 4'h0;
assign TX_DATA_34_const_net_0              = 4'h0;
assign TX_DATA_35_const_net_0              = 4'h0;
assign TX_DATA_36_const_net_0              = 4'h0;
assign TX_DATA_37_const_net_0              = 4'h0;
assign TX_DATA_38_const_net_0              = 4'h0;
assign TX_DATA_39_const_net_0              = 4'h0;
assign TX_DATA_40_const_net_0              = 4'h0;
assign TX_DATA_41_const_net_0              = 4'h0;
assign TX_DATA_42_const_net_0              = 4'h0;
assign TX_DATA_43_const_net_0              = 4'h0;
assign TX_DATA_44_const_net_0              = 4'h0;
assign TX_DATA_45_const_net_0              = 4'h0;
assign TX_DATA_46_const_net_0              = 4'h0;
assign TX_DATA_47_const_net_0              = 4'h0;
assign TX_DATA_48_const_net_0              = 4'h0;
assign TX_DATA_49_const_net_0              = 4'h0;
assign TX_DATA_50_const_net_0              = 4'h0;
assign TX_DATA_51_const_net_0              = 4'h0;
assign TX_DATA_52_const_net_0              = 4'h0;
assign TX_DATA_53_const_net_0              = 4'h0;
assign TX_DATA_54_const_net_0              = 4'h0;
assign TX_DATA_55_const_net_0              = 4'h0;
assign TX_DATA_56_const_net_0              = 4'h0;
assign TX_DATA_57_const_net_0              = 4'h0;
assign TX_DATA_58_const_net_0              = 4'h0;
assign TX_DATA_59_const_net_0              = 4'h0;
assign TX_DATA_60_const_net_0              = 4'h0;
assign TX_DATA_61_const_net_0              = 4'h0;
assign TX_DATA_62_const_net_0              = 4'h0;
assign TX_DATA_63_const_net_0              = 4'h0;
assign TX_DATA_64_const_net_0              = 4'h0;
assign TX_DATA_65_const_net_0              = 4'h0;
assign TX_DATA_66_const_net_0              = 4'h0;
assign TX_DATA_67_const_net_0              = 4'h0;
assign TX_DATA_68_const_net_0              = 4'h0;
assign TX_DATA_69_const_net_0              = 4'h0;
assign TX_DATA_70_const_net_0              = 4'h0;
assign TX_DATA_71_const_net_0              = 4'h0;
assign TX_DATA_72_const_net_0              = 4'h0;
assign TX_DATA_73_const_net_0              = 4'h0;
assign TX_DATA_74_const_net_0              = 4'h0;
assign TX_DATA_75_const_net_0              = 4'h0;
assign TX_DATA_76_const_net_0              = 4'h0;
assign TX_DATA_77_const_net_0              = 4'h0;
assign TX_DATA_78_const_net_0              = 4'h0;
assign TX_DATA_79_const_net_0              = 4'h0;
assign TX_DATA_80_const_net_0              = 4'h0;
assign TX_DATA_81_const_net_0              = 4'h0;
assign TX_DATA_82_const_net_0              = 4'h0;
assign TX_DATA_83_const_net_0              = 4'h0;
assign TX_DATA_84_const_net_0              = 4'h0;
assign TX_DATA_85_const_net_0              = 4'h0;
assign TX_DATA_86_const_net_0              = 4'h0;
assign TX_DATA_87_const_net_0              = 4'h0;
assign TX_DATA_88_const_net_0              = 4'h0;
assign TX_DATA_89_const_net_0              = 4'h0;
assign TX_DATA_90_const_net_0              = 4'h0;
assign TX_DATA_91_const_net_0              = 4'h0;
assign TX_DATA_92_const_net_0              = 4'h0;
assign TX_DATA_93_const_net_0              = 4'h0;
assign TX_DATA_94_const_net_0              = 4'h0;
assign TX_DATA_95_const_net_0              = 4'h0;
assign TX_DATA_96_const_net_0              = 4'h0;
assign TX_DATA_97_const_net_0              = 4'h0;
assign TX_DATA_98_const_net_0              = 4'h0;
assign TX_DATA_99_const_net_0              = 4'h0;
assign TX_DATA_100_const_net_0             = 4'h0;
assign TX_DATA_101_const_net_0             = 4'h0;
assign TX_DATA_102_const_net_0             = 4'h0;
assign TX_DATA_103_const_net_0             = 4'h0;
assign TX_DATA_104_const_net_0             = 4'h0;
assign TX_DATA_105_const_net_0             = 4'h0;
assign TX_DATA_106_const_net_0             = 4'h0;
assign TX_DATA_107_const_net_0             = 4'h0;
assign TX_DATA_108_const_net_0             = 4'h0;
assign TX_DATA_109_const_net_0             = 4'h0;
assign TX_DATA_110_const_net_0             = 4'h0;
assign TX_DATA_111_const_net_0             = 4'h0;
assign TX_DATA_112_const_net_0             = 4'h0;
assign TX_DATA_113_const_net_0             = 4'h0;
assign TX_DATA_114_const_net_0             = 4'h0;
assign TX_DATA_115_const_net_0             = 4'h0;
assign TX_DATA_116_const_net_0             = 4'h0;
assign TX_DATA_117_const_net_0             = 4'h0;
assign TX_DATA_118_const_net_0             = 4'h0;
assign TX_DATA_119_const_net_0             = 4'h0;
assign TX_DATA_120_const_net_0             = 4'h0;
assign TX_DATA_121_const_net_0             = 4'h0;
assign TX_DATA_122_const_net_0             = 4'h0;
assign TX_DATA_123_const_net_0             = 4'h0;
assign TX_DATA_124_const_net_0             = 4'h0;
assign TX_DATA_125_const_net_0             = 4'h0;
assign TX_DATA_126_const_net_0             = 4'h0;
assign TX_DATA_127_const_net_0             = 4'h0;
assign OE_DATA_12_const_net_0              = 4'h0;
assign OE_DATA_13_const_net_0              = 4'h0;
assign OE_DATA_14_const_net_0              = 4'h0;
assign OE_DATA_15_const_net_0              = 4'h0;
assign OE_DATA_16_const_net_0              = 4'h0;
assign OE_DATA_17_const_net_0              = 4'h0;
assign OE_DATA_18_const_net_0              = 4'h0;
assign OE_DATA_19_const_net_0              = 4'h0;
assign OE_DATA_20_const_net_0              = 4'h0;
assign OE_DATA_21_const_net_0              = 4'h0;
assign OE_DATA_22_const_net_0              = 4'h0;
assign OE_DATA_23_const_net_0              = 4'h0;
assign OE_DATA_24_const_net_0              = 4'h0;
assign OE_DATA_25_const_net_0              = 4'h0;
assign OE_DATA_26_const_net_0              = 4'h0;
assign OE_DATA_27_const_net_0              = 4'h0;
assign OE_DATA_28_const_net_0              = 4'h0;
assign OE_DATA_29_const_net_0              = 4'h0;
assign OE_DATA_30_const_net_0              = 4'h0;
assign OE_DATA_31_const_net_0              = 4'h0;
assign OE_DATA_32_const_net_0              = 4'h0;
assign OE_DATA_33_const_net_0              = 4'h0;
assign OE_DATA_34_const_net_0              = 4'h0;
assign OE_DATA_35_const_net_0              = 4'h0;
assign OE_DATA_36_const_net_0              = 4'h0;
assign OE_DATA_37_const_net_0              = 4'h0;
assign OE_DATA_38_const_net_0              = 4'h0;
assign OE_DATA_39_const_net_0              = 4'h0;
assign OE_DATA_40_const_net_0              = 4'h0;
assign OE_DATA_41_const_net_0              = 4'h0;
assign OE_DATA_42_const_net_0              = 4'h0;
assign OE_DATA_43_const_net_0              = 4'h0;
assign OE_DATA_44_const_net_0              = 4'h0;
assign OE_DATA_45_const_net_0              = 4'h0;
assign OE_DATA_46_const_net_0              = 4'h0;
assign OE_DATA_47_const_net_0              = 4'h0;
assign OE_DATA_48_const_net_0              = 4'h0;
assign OE_DATA_49_const_net_0              = 4'h0;
assign OE_DATA_50_const_net_0              = 4'h0;
assign OE_DATA_51_const_net_0              = 4'h0;
assign OE_DATA_52_const_net_0              = 4'h0;
assign OE_DATA_53_const_net_0              = 4'h0;
assign OE_DATA_54_const_net_0              = 4'h0;
assign OE_DATA_55_const_net_0              = 4'h0;
assign OE_DATA_56_const_net_0              = 4'h0;
assign OE_DATA_57_const_net_0              = 4'h0;
assign OE_DATA_58_const_net_0              = 4'h0;
assign OE_DATA_59_const_net_0              = 4'h0;
assign OE_DATA_60_const_net_0              = 4'h0;
assign OE_DATA_61_const_net_0              = 4'h0;
assign OE_DATA_62_const_net_0              = 4'h0;
assign OE_DATA_63_const_net_0              = 4'h0;
assign OE_DATA_64_const_net_0              = 4'h0;
assign OE_DATA_65_const_net_0              = 4'h0;
assign OE_DATA_66_const_net_0              = 4'h0;
assign OE_DATA_67_const_net_0              = 4'h0;
assign OE_DATA_68_const_net_0              = 4'h0;
assign OE_DATA_69_const_net_0              = 4'h0;
assign OE_DATA_70_const_net_0              = 4'h0;
assign OE_DATA_71_const_net_0              = 4'h0;
assign OE_DATA_72_const_net_0              = 4'h0;
assign OE_DATA_73_const_net_0              = 4'h0;
assign OE_DATA_74_const_net_0              = 4'h0;
assign OE_DATA_75_const_net_0              = 4'h0;
assign OE_DATA_76_const_net_0              = 4'h0;
assign OE_DATA_77_const_net_0              = 4'h0;
assign OE_DATA_78_const_net_0              = 4'h0;
assign OE_DATA_79_const_net_0              = 4'h0;
assign OE_DATA_80_const_net_0              = 4'h0;
assign OE_DATA_81_const_net_0              = 4'h0;
assign OE_DATA_82_const_net_0              = 4'h0;
assign OE_DATA_83_const_net_0              = 4'h0;
assign OE_DATA_84_const_net_0              = 4'h0;
assign OE_DATA_85_const_net_0              = 4'h0;
assign OE_DATA_86_const_net_0              = 4'h0;
assign OE_DATA_87_const_net_0              = 4'h0;
assign OE_DATA_88_const_net_0              = 4'h0;
assign OE_DATA_89_const_net_0              = 4'h0;
assign OE_DATA_90_const_net_0              = 4'h0;
assign OE_DATA_91_const_net_0              = 4'h0;
assign OE_DATA_92_const_net_0              = 4'h0;
assign OE_DATA_93_const_net_0              = 4'h0;
assign OE_DATA_94_const_net_0              = 4'h0;
assign OE_DATA_95_const_net_0              = 4'h0;
assign OE_DATA_96_const_net_0              = 4'h0;
assign OE_DATA_97_const_net_0              = 4'h0;
assign OE_DATA_98_const_net_0              = 4'h0;
assign OE_DATA_99_const_net_0              = 4'h0;
assign OE_DATA_100_const_net_0             = 4'h0;
assign OE_DATA_101_const_net_0             = 4'h0;
assign OE_DATA_102_const_net_0             = 4'h0;
assign OE_DATA_103_const_net_0             = 4'h0;
assign OE_DATA_104_const_net_0             = 4'h0;
assign OE_DATA_105_const_net_0             = 4'h0;
assign OE_DATA_106_const_net_0             = 4'h0;
assign OE_DATA_107_const_net_0             = 4'h0;
assign OE_DATA_108_const_net_0             = 4'h0;
assign OE_DATA_109_const_net_0             = 4'h0;
assign OE_DATA_110_const_net_0             = 4'h0;
assign OE_DATA_111_const_net_0             = 4'h0;
assign OE_DATA_112_const_net_0             = 4'h0;
assign OE_DATA_113_const_net_0             = 4'h0;
assign OE_DATA_114_const_net_0             = 4'h0;
assign OE_DATA_115_const_net_0             = 4'h0;
assign OE_DATA_116_const_net_0             = 4'h0;
assign OE_DATA_117_const_net_0             = 4'h0;
assign OE_DATA_118_const_net_0             = 4'h0;
assign OE_DATA_119_const_net_0             = 4'h0;
assign OE_DATA_120_const_net_0             = 4'h0;
assign OE_DATA_121_const_net_0             = 4'h0;
assign OE_DATA_122_const_net_0             = 4'h0;
assign OE_DATA_123_const_net_0             = 4'h0;
assign OE_DATA_124_const_net_0             = 4'h0;
assign OE_DATA_125_const_net_0             = 4'h0;
assign OE_DATA_126_const_net_0             = 4'h0;
assign OE_DATA_127_const_net_0             = 4'h0;
assign PAD_const_net_0                     = 12'h000;
assign PAD_I_const_net_0                   = 12'h000;
assign PAD_N_const_net_0                   = 12'h000;
assign PAD_I_N_const_net_0                 = 12'h000;
assign RX_DQS_90_const_net_1               = 2'h0;
assign FIFO_WR_PTR_const_net_1             = 3'h0;
assign FIFO_RD_PTR_const_net_1             = 3'h0;
assign EYE_MONITOR_LANE_WIDTH_const_net_1  = 3'h0;
assign TX_DATA_1_const_net_0               = 4'h0;
assign TX_DATA_2_const_net_0               = 4'h0;
assign TX_DATA_3_const_net_0               = 4'h0;
assign TX_DATA_4_const_net_0               = 4'h0;
assign TX_DATA_5_const_net_0               = 4'h0;
assign TX_DATA_6_const_net_0               = 4'h0;
assign TX_DATA_7_const_net_0               = 4'h0;
assign TX_DATA_8_const_net_0               = 4'h0;
assign TX_DATA_9_const_net_0               = 4'h0;
assign TX_DATA_10_const_net_0              = 4'h0;
assign TX_DATA_11_const_net_0              = 4'h0;
assign TX_DATA_12_const_net_1              = 4'h0;
assign TX_DATA_13_const_net_1              = 4'h0;
assign TX_DATA_14_const_net_1              = 4'h0;
assign TX_DATA_15_const_net_1              = 4'h0;
assign TX_DATA_16_const_net_1              = 4'h0;
assign TX_DATA_17_const_net_1              = 4'h0;
assign TX_DATA_18_const_net_1              = 4'h0;
assign TX_DATA_19_const_net_1              = 4'h0;
assign TX_DATA_20_const_net_1              = 4'h0;
assign TX_DATA_21_const_net_1              = 4'h0;
assign TX_DATA_22_const_net_1              = 4'h0;
assign TX_DATA_23_const_net_1              = 4'h0;
assign TX_DATA_24_const_net_1              = 4'h0;
assign TX_DATA_25_const_net_1              = 4'h0;
assign TX_DATA_26_const_net_1              = 4'h0;
assign TX_DATA_27_const_net_1              = 4'h0;
assign TX_DATA_28_const_net_1              = 4'h0;
assign TX_DATA_29_const_net_1              = 4'h0;
assign TX_DATA_30_const_net_1              = 4'h0;
assign TX_DATA_31_const_net_1              = 4'h0;
assign TX_DATA_32_const_net_1              = 4'h0;
assign TX_DATA_33_const_net_1              = 4'h0;
assign TX_DATA_34_const_net_1              = 4'h0;
assign TX_DATA_35_const_net_1              = 4'h0;
assign TX_DATA_36_const_net_1              = 4'h0;
assign TX_DATA_37_const_net_1              = 4'h0;
assign TX_DATA_38_const_net_1              = 4'h0;
assign TX_DATA_39_const_net_1              = 4'h0;
assign TX_DATA_40_const_net_1              = 4'h0;
assign TX_DATA_41_const_net_1              = 4'h0;
assign TX_DATA_42_const_net_1              = 4'h0;
assign TX_DATA_43_const_net_1              = 4'h0;
assign TX_DATA_44_const_net_1              = 4'h0;
assign TX_DATA_45_const_net_1              = 4'h0;
assign TX_DATA_46_const_net_1              = 4'h0;
assign TX_DATA_47_const_net_1              = 4'h0;
assign TX_DATA_48_const_net_1              = 4'h0;
assign TX_DATA_49_const_net_1              = 4'h0;
assign TX_DATA_50_const_net_1              = 4'h0;
assign TX_DATA_51_const_net_1              = 4'h0;
assign TX_DATA_52_const_net_1              = 4'h0;
assign TX_DATA_53_const_net_1              = 4'h0;
assign TX_DATA_54_const_net_1              = 4'h0;
assign TX_DATA_55_const_net_1              = 4'h0;
assign TX_DATA_56_const_net_1              = 4'h0;
assign TX_DATA_57_const_net_1              = 4'h0;
assign TX_DATA_58_const_net_1              = 4'h0;
assign TX_DATA_59_const_net_1              = 4'h0;
assign TX_DATA_60_const_net_1              = 4'h0;
assign TX_DATA_61_const_net_1              = 4'h0;
assign TX_DATA_62_const_net_1              = 4'h0;
assign TX_DATA_63_const_net_1              = 4'h0;
assign TX_DATA_64_const_net_1              = 4'h0;
assign TX_DATA_65_const_net_1              = 4'h0;
assign TX_DATA_66_const_net_1              = 4'h0;
assign TX_DATA_67_const_net_1              = 4'h0;
assign TX_DATA_68_const_net_1              = 4'h0;
assign TX_DATA_69_const_net_1              = 4'h0;
assign TX_DATA_70_const_net_1              = 4'h0;
assign TX_DATA_71_const_net_1              = 4'h0;
assign TX_DATA_72_const_net_1              = 4'h0;
assign TX_DATA_73_const_net_1              = 4'h0;
assign TX_DATA_74_const_net_1              = 4'h0;
assign TX_DATA_75_const_net_1              = 4'h0;
assign TX_DATA_76_const_net_1              = 4'h0;
assign TX_DATA_77_const_net_1              = 4'h0;
assign TX_DATA_78_const_net_1              = 4'h0;
assign TX_DATA_79_const_net_1              = 4'h0;
assign TX_DATA_80_const_net_1              = 4'h0;
assign TX_DATA_81_const_net_1              = 4'h0;
assign TX_DATA_82_const_net_1              = 4'h0;
assign TX_DATA_83_const_net_1              = 4'h0;
assign TX_DATA_84_const_net_1              = 4'h0;
assign TX_DATA_85_const_net_1              = 4'h0;
assign TX_DATA_86_const_net_1              = 4'h0;
assign TX_DATA_87_const_net_1              = 4'h0;
assign TX_DATA_88_const_net_1              = 4'h0;
assign TX_DATA_89_const_net_1              = 4'h0;
assign TX_DATA_90_const_net_1              = 4'h0;
assign TX_DATA_91_const_net_1              = 4'h0;
assign TX_DATA_92_const_net_1              = 4'h0;
assign TX_DATA_93_const_net_1              = 4'h0;
assign TX_DATA_94_const_net_1              = 4'h0;
assign TX_DATA_95_const_net_1              = 4'h0;
assign TX_DATA_96_const_net_1              = 4'h0;
assign TX_DATA_97_const_net_1              = 4'h0;
assign TX_DATA_98_const_net_1              = 4'h0;
assign TX_DATA_99_const_net_1              = 4'h0;
assign TX_DATA_100_const_net_1             = 4'h0;
assign TX_DATA_101_const_net_1             = 4'h0;
assign TX_DATA_102_const_net_1             = 4'h0;
assign TX_DATA_103_const_net_1             = 4'h0;
assign TX_DATA_104_const_net_1             = 4'h0;
assign TX_DATA_105_const_net_1             = 4'h0;
assign TX_DATA_106_const_net_1             = 4'h0;
assign TX_DATA_107_const_net_1             = 4'h0;
assign TX_DATA_108_const_net_1             = 4'h0;
assign TX_DATA_109_const_net_1             = 4'h0;
assign TX_DATA_110_const_net_1             = 4'h0;
assign TX_DATA_111_const_net_1             = 4'h0;
assign TX_DATA_112_const_net_1             = 4'h0;
assign TX_DATA_113_const_net_1             = 4'h0;
assign TX_DATA_114_const_net_1             = 4'h0;
assign TX_DATA_115_const_net_1             = 4'h0;
assign TX_DATA_116_const_net_1             = 4'h0;
assign TX_DATA_117_const_net_1             = 4'h0;
assign TX_DATA_118_const_net_1             = 4'h0;
assign TX_DATA_119_const_net_1             = 4'h0;
assign TX_DATA_120_const_net_1             = 4'h0;
assign TX_DATA_121_const_net_1             = 4'h0;
assign TX_DATA_122_const_net_1             = 4'h0;
assign TX_DATA_123_const_net_1             = 4'h0;
assign TX_DATA_124_const_net_1             = 4'h0;
assign TX_DATA_125_const_net_1             = 4'h0;
assign TX_DATA_126_const_net_1             = 4'h0;
assign TX_DATA_127_const_net_1             = 4'h0;
assign OE_DATA_1_const_net_3               = 4'h0;
assign OE_DATA_2_const_net_1               = 4'h0;
assign OE_DATA_3_const_net_1               = 4'h0;
assign OE_DATA_4_const_net_1               = 4'h0;
assign OE_DATA_5_const_net_1               = 4'h0;
assign OE_DATA_6_const_net_1               = 4'h0;
assign OE_DATA_7_const_net_1               = 4'h0;
assign OE_DATA_8_const_net_1               = 4'h0;
assign OE_DATA_9_const_net_1               = 4'h0;
assign OE_DATA_10_const_net_1              = 4'h0;
assign OE_DATA_11_const_net_1              = 4'h0;
assign OE_DATA_12_const_net_1              = 4'h0;
assign OE_DATA_13_const_net_1              = 4'h0;
assign OE_DATA_14_const_net_1              = 4'h0;
assign OE_DATA_15_const_net_1              = 4'h0;
assign OE_DATA_16_const_net_1              = 4'h0;
assign OE_DATA_17_const_net_1              = 4'h0;
assign OE_DATA_18_const_net_1              = 4'h0;
assign OE_DATA_19_const_net_1              = 4'h0;
assign OE_DATA_20_const_net_1              = 4'h0;
assign OE_DATA_21_const_net_1              = 4'h0;
assign OE_DATA_22_const_net_1              = 4'h0;
assign OE_DATA_23_const_net_1              = 4'h0;
assign OE_DATA_24_const_net_1              = 4'h0;
assign OE_DATA_25_const_net_1              = 4'h0;
assign OE_DATA_26_const_net_1              = 4'h0;
assign OE_DATA_27_const_net_1              = 4'h0;
assign OE_DATA_28_const_net_1              = 4'h0;
assign OE_DATA_29_const_net_1              = 4'h0;
assign OE_DATA_30_const_net_1              = 4'h0;
assign OE_DATA_31_const_net_1              = 4'h0;
assign OE_DATA_32_const_net_1              = 4'h0;
assign OE_DATA_33_const_net_1              = 4'h0;
assign OE_DATA_34_const_net_1              = 4'h0;
assign OE_DATA_35_const_net_1              = 4'h0;
assign OE_DATA_36_const_net_1              = 4'h0;
assign OE_DATA_37_const_net_1              = 4'h0;
assign OE_DATA_38_const_net_1              = 4'h0;
assign OE_DATA_39_const_net_1              = 4'h0;
assign OE_DATA_40_const_net_1              = 4'h0;
assign OE_DATA_41_const_net_1              = 4'h0;
assign OE_DATA_42_const_net_1              = 4'h0;
assign OE_DATA_43_const_net_1              = 4'h0;
assign OE_DATA_44_const_net_1              = 4'h0;
assign OE_DATA_45_const_net_1              = 4'h0;
assign OE_DATA_46_const_net_1              = 4'h0;
assign OE_DATA_47_const_net_1              = 4'h0;
assign OE_DATA_48_const_net_1              = 4'h0;
assign OE_DATA_49_const_net_1              = 4'h0;
assign OE_DATA_50_const_net_1              = 4'h0;
assign OE_DATA_51_const_net_1              = 4'h0;
assign OE_DATA_52_const_net_1              = 4'h0;
assign OE_DATA_53_const_net_1              = 4'h0;
assign OE_DATA_54_const_net_1              = 4'h0;
assign OE_DATA_55_const_net_1              = 4'h0;
assign OE_DATA_56_const_net_1              = 4'h0;
assign OE_DATA_57_const_net_1              = 4'h0;
assign OE_DATA_58_const_net_1              = 4'h0;
assign OE_DATA_59_const_net_1              = 4'h0;
assign OE_DATA_60_const_net_1              = 4'h0;
assign OE_DATA_61_const_net_1              = 4'h0;
assign OE_DATA_62_const_net_1              = 4'h0;
assign OE_DATA_63_const_net_1              = 4'h0;
assign OE_DATA_64_const_net_1              = 4'h0;
assign OE_DATA_65_const_net_1              = 4'h0;
assign OE_DATA_66_const_net_1              = 4'h0;
assign OE_DATA_67_const_net_1              = 4'h0;
assign OE_DATA_68_const_net_1              = 4'h0;
assign OE_DATA_69_const_net_1              = 4'h0;
assign OE_DATA_70_const_net_1              = 4'h0;
assign OE_DATA_71_const_net_1              = 4'h0;
assign OE_DATA_72_const_net_1              = 4'h0;
assign OE_DATA_73_const_net_1              = 4'h0;
assign OE_DATA_74_const_net_1              = 4'h0;
assign OE_DATA_75_const_net_1              = 4'h0;
assign OE_DATA_76_const_net_1              = 4'h0;
assign OE_DATA_77_const_net_1              = 4'h0;
assign OE_DATA_78_const_net_1              = 4'h0;
assign OE_DATA_79_const_net_1              = 4'h0;
assign OE_DATA_80_const_net_1              = 4'h0;
assign OE_DATA_81_const_net_1              = 4'h0;
assign OE_DATA_82_const_net_1              = 4'h0;
assign OE_DATA_83_const_net_1              = 4'h0;
assign OE_DATA_84_const_net_1              = 4'h0;
assign OE_DATA_85_const_net_1              = 4'h0;
assign OE_DATA_86_const_net_1              = 4'h0;
assign OE_DATA_87_const_net_1              = 4'h0;
assign OE_DATA_88_const_net_1              = 4'h0;
assign OE_DATA_89_const_net_1              = 4'h0;
assign OE_DATA_90_const_net_1              = 4'h0;
assign OE_DATA_91_const_net_1              = 4'h0;
assign OE_DATA_92_const_net_1              = 4'h0;
assign OE_DATA_93_const_net_1              = 4'h0;
assign OE_DATA_94_const_net_1              = 4'h0;
assign OE_DATA_95_const_net_1              = 4'h0;
assign OE_DATA_96_const_net_1              = 4'h0;
assign OE_DATA_97_const_net_1              = 4'h0;
assign OE_DATA_98_const_net_1              = 4'h0;
assign OE_DATA_99_const_net_1              = 4'h0;
assign OE_DATA_100_const_net_1             = 4'h0;
assign OE_DATA_101_const_net_1             = 4'h0;
assign OE_DATA_102_const_net_1             = 4'h0;
assign OE_DATA_103_const_net_1             = 4'h0;
assign OE_DATA_104_const_net_1             = 4'h0;
assign OE_DATA_105_const_net_1             = 4'h0;
assign OE_DATA_106_const_net_1             = 4'h0;
assign OE_DATA_107_const_net_1             = 4'h0;
assign OE_DATA_108_const_net_1             = 4'h0;
assign OE_DATA_109_const_net_1             = 4'h0;
assign OE_DATA_110_const_net_1             = 4'h0;
assign OE_DATA_111_const_net_1             = 4'h0;
assign OE_DATA_112_const_net_1             = 4'h0;
assign OE_DATA_113_const_net_1             = 4'h0;
assign OE_DATA_114_const_net_1             = 4'h0;
assign OE_DATA_115_const_net_1             = 4'h0;
assign OE_DATA_116_const_net_1             = 4'h0;
assign OE_DATA_117_const_net_1             = 4'h0;
assign OE_DATA_118_const_net_1             = 4'h0;
assign OE_DATA_119_const_net_1             = 4'h0;
assign OE_DATA_120_const_net_1             = 4'h0;
assign OE_DATA_121_const_net_1             = 4'h0;
assign OE_DATA_122_const_net_1             = 4'h0;
assign OE_DATA_123_const_net_1             = 4'h0;
assign OE_DATA_124_const_net_1             = 4'h0;
assign OE_DATA_125_const_net_1             = 4'h0;
assign OE_DATA_126_const_net_1             = 4'h0;
assign OE_DATA_127_const_net_1             = 4'h0;
assign RX_DQS_90_const_net_2               = 2'h0;
assign FIFO_WR_PTR_const_net_2             = 3'h0;
assign FIFO_RD_PTR_const_net_2             = 3'h0;
assign EYE_MONITOR_LANE_WIDTH_const_net_2  = 3'h0;
assign TX_DATA_1_const_net_1               = 4'h0;
assign TX_DATA_2_const_net_1               = 4'h0;
assign TX_DATA_3_const_net_1               = 4'h0;
assign TX_DATA_4_const_net_1               = 4'h0;
assign TX_DATA_5_const_net_1               = 4'h0;
assign TX_DATA_6_const_net_1               = 4'h0;
assign TX_DATA_7_const_net_1               = 4'h0;
assign TX_DATA_8_const_net_1               = 4'h0;
assign TX_DATA_9_const_net_1               = 4'h0;
assign TX_DATA_10_const_net_1              = 4'h0;
assign TX_DATA_11_const_net_1              = 4'h0;
assign TX_DATA_12_const_net_2              = 4'h0;
assign TX_DATA_13_const_net_2              = 4'h0;
assign TX_DATA_14_const_net_2              = 4'h0;
assign TX_DATA_15_const_net_2              = 4'h0;
assign TX_DATA_16_const_net_2              = 4'h0;
assign TX_DATA_17_const_net_2              = 4'h0;
assign TX_DATA_18_const_net_2              = 4'h0;
assign TX_DATA_19_const_net_2              = 4'h0;
assign TX_DATA_20_const_net_2              = 4'h0;
assign TX_DATA_21_const_net_2              = 4'h0;
assign TX_DATA_22_const_net_2              = 4'h0;
assign TX_DATA_23_const_net_2              = 4'h0;
assign TX_DATA_24_const_net_2              = 4'h0;
assign TX_DATA_25_const_net_2              = 4'h0;
assign TX_DATA_26_const_net_2              = 4'h0;
assign TX_DATA_27_const_net_2              = 4'h0;
assign TX_DATA_28_const_net_2              = 4'h0;
assign TX_DATA_29_const_net_2              = 4'h0;
assign TX_DATA_30_const_net_2              = 4'h0;
assign TX_DATA_31_const_net_2              = 4'h0;
assign TX_DATA_32_const_net_2              = 4'h0;
assign TX_DATA_33_const_net_2              = 4'h0;
assign TX_DATA_34_const_net_2              = 4'h0;
assign TX_DATA_35_const_net_2              = 4'h0;
assign TX_DATA_36_const_net_2              = 4'h0;
assign TX_DATA_37_const_net_2              = 4'h0;
assign TX_DATA_38_const_net_2              = 4'h0;
assign TX_DATA_39_const_net_2              = 4'h0;
assign TX_DATA_40_const_net_2              = 4'h0;
assign TX_DATA_41_const_net_2              = 4'h0;
assign TX_DATA_42_const_net_2              = 4'h0;
assign TX_DATA_43_const_net_2              = 4'h0;
assign TX_DATA_44_const_net_2              = 4'h0;
assign TX_DATA_45_const_net_2              = 4'h0;
assign TX_DATA_46_const_net_2              = 4'h0;
assign TX_DATA_47_const_net_2              = 4'h0;
assign TX_DATA_48_const_net_2              = 4'h0;
assign TX_DATA_49_const_net_2              = 4'h0;
assign TX_DATA_50_const_net_2              = 4'h0;
assign TX_DATA_51_const_net_2              = 4'h0;
assign TX_DATA_52_const_net_2              = 4'h0;
assign TX_DATA_53_const_net_2              = 4'h0;
assign TX_DATA_54_const_net_2              = 4'h0;
assign TX_DATA_55_const_net_2              = 4'h0;
assign TX_DATA_56_const_net_2              = 4'h0;
assign TX_DATA_57_const_net_2              = 4'h0;
assign TX_DATA_58_const_net_2              = 4'h0;
assign TX_DATA_59_const_net_2              = 4'h0;
assign TX_DATA_60_const_net_2              = 4'h0;
assign TX_DATA_61_const_net_2              = 4'h0;
assign TX_DATA_62_const_net_2              = 4'h0;
assign TX_DATA_63_const_net_2              = 4'h0;
assign TX_DATA_64_const_net_2              = 4'h0;
assign TX_DATA_65_const_net_2              = 4'h0;
assign TX_DATA_66_const_net_2              = 4'h0;
assign TX_DATA_67_const_net_2              = 4'h0;
assign TX_DATA_68_const_net_2              = 4'h0;
assign TX_DATA_69_const_net_2              = 4'h0;
assign TX_DATA_70_const_net_2              = 4'h0;
assign TX_DATA_71_const_net_2              = 4'h0;
assign TX_DATA_72_const_net_2              = 4'h0;
assign TX_DATA_73_const_net_2              = 4'h0;
assign TX_DATA_74_const_net_2              = 4'h0;
assign TX_DATA_75_const_net_2              = 4'h0;
assign TX_DATA_76_const_net_2              = 4'h0;
assign TX_DATA_77_const_net_2              = 4'h0;
assign TX_DATA_78_const_net_2              = 4'h0;
assign TX_DATA_79_const_net_2              = 4'h0;
assign TX_DATA_80_const_net_2              = 4'h0;
assign TX_DATA_81_const_net_2              = 4'h0;
assign TX_DATA_82_const_net_2              = 4'h0;
assign TX_DATA_83_const_net_2              = 4'h0;
assign TX_DATA_84_const_net_2              = 4'h0;
assign TX_DATA_85_const_net_2              = 4'h0;
assign TX_DATA_86_const_net_2              = 4'h0;
assign TX_DATA_87_const_net_2              = 4'h0;
assign TX_DATA_88_const_net_2              = 4'h0;
assign TX_DATA_89_const_net_2              = 4'h0;
assign TX_DATA_90_const_net_2              = 4'h0;
assign TX_DATA_91_const_net_2              = 4'h0;
assign TX_DATA_92_const_net_2              = 4'h0;
assign TX_DATA_93_const_net_2              = 4'h0;
assign TX_DATA_94_const_net_2              = 4'h0;
assign TX_DATA_95_const_net_2              = 4'h0;
assign TX_DATA_96_const_net_2              = 4'h0;
assign TX_DATA_97_const_net_2              = 4'h0;
assign TX_DATA_98_const_net_2              = 4'h0;
assign TX_DATA_99_const_net_2              = 4'h0;
assign TX_DATA_100_const_net_2             = 4'h0;
assign TX_DATA_101_const_net_2             = 4'h0;
assign TX_DATA_102_const_net_2             = 4'h0;
assign TX_DATA_103_const_net_2             = 4'h0;
assign TX_DATA_104_const_net_2             = 4'h0;
assign TX_DATA_105_const_net_2             = 4'h0;
assign TX_DATA_106_const_net_2             = 4'h0;
assign TX_DATA_107_const_net_2             = 4'h0;
assign TX_DATA_108_const_net_2             = 4'h0;
assign TX_DATA_109_const_net_2             = 4'h0;
assign TX_DATA_110_const_net_2             = 4'h0;
assign TX_DATA_111_const_net_2             = 4'h0;
assign TX_DATA_112_const_net_2             = 4'h0;
assign TX_DATA_113_const_net_2             = 4'h0;
assign TX_DATA_114_const_net_2             = 4'h0;
assign TX_DATA_115_const_net_2             = 4'h0;
assign TX_DATA_116_const_net_2             = 4'h0;
assign TX_DATA_117_const_net_2             = 4'h0;
assign TX_DATA_118_const_net_2             = 4'h0;
assign TX_DATA_119_const_net_2             = 4'h0;
assign TX_DATA_120_const_net_2             = 4'h0;
assign TX_DATA_121_const_net_2             = 4'h0;
assign TX_DATA_122_const_net_2             = 4'h0;
assign TX_DATA_123_const_net_2             = 4'h0;
assign TX_DATA_124_const_net_2             = 4'h0;
assign TX_DATA_125_const_net_2             = 4'h0;
assign TX_DATA_126_const_net_2             = 4'h0;
assign TX_DATA_127_const_net_2             = 4'h0;
assign OE_DATA_1_const_net_4               = 4'h0;
assign OE_DATA_2_const_net_2               = 4'h0;
assign OE_DATA_3_const_net_2               = 4'h0;
assign OE_DATA_4_const_net_2               = 4'h0;
assign OE_DATA_5_const_net_2               = 4'h0;
assign OE_DATA_6_const_net_2               = 4'h0;
assign OE_DATA_7_const_net_2               = 4'h0;
assign OE_DATA_8_const_net_2               = 4'h0;
assign OE_DATA_9_const_net_2               = 4'h0;
assign OE_DATA_10_const_net_2              = 4'h0;
assign OE_DATA_11_const_net_2              = 4'h0;
assign OE_DATA_12_const_net_2              = 4'h0;
assign OE_DATA_13_const_net_2              = 4'h0;
assign OE_DATA_14_const_net_2              = 4'h0;
assign OE_DATA_15_const_net_2              = 4'h0;
assign OE_DATA_16_const_net_2              = 4'h0;
assign OE_DATA_17_const_net_2              = 4'h0;
assign OE_DATA_18_const_net_2              = 4'h0;
assign OE_DATA_19_const_net_2              = 4'h0;
assign OE_DATA_20_const_net_2              = 4'h0;
assign OE_DATA_21_const_net_2              = 4'h0;
assign OE_DATA_22_const_net_2              = 4'h0;
assign OE_DATA_23_const_net_2              = 4'h0;
assign OE_DATA_24_const_net_2              = 4'h0;
assign OE_DATA_25_const_net_2              = 4'h0;
assign OE_DATA_26_const_net_2              = 4'h0;
assign OE_DATA_27_const_net_2              = 4'h0;
assign OE_DATA_28_const_net_2              = 4'h0;
assign OE_DATA_29_const_net_2              = 4'h0;
assign OE_DATA_30_const_net_2              = 4'h0;
assign OE_DATA_31_const_net_2              = 4'h0;
assign OE_DATA_32_const_net_2              = 4'h0;
assign OE_DATA_33_const_net_2              = 4'h0;
assign OE_DATA_34_const_net_2              = 4'h0;
assign OE_DATA_35_const_net_2              = 4'h0;
assign OE_DATA_36_const_net_2              = 4'h0;
assign OE_DATA_37_const_net_2              = 4'h0;
assign OE_DATA_38_const_net_2              = 4'h0;
assign OE_DATA_39_const_net_2              = 4'h0;
assign OE_DATA_40_const_net_2              = 4'h0;
assign OE_DATA_41_const_net_2              = 4'h0;
assign OE_DATA_42_const_net_2              = 4'h0;
assign OE_DATA_43_const_net_2              = 4'h0;
assign OE_DATA_44_const_net_2              = 4'h0;
assign OE_DATA_45_const_net_2              = 4'h0;
assign OE_DATA_46_const_net_2              = 4'h0;
assign OE_DATA_47_const_net_2              = 4'h0;
assign OE_DATA_48_const_net_2              = 4'h0;
assign OE_DATA_49_const_net_2              = 4'h0;
assign OE_DATA_50_const_net_2              = 4'h0;
assign OE_DATA_51_const_net_2              = 4'h0;
assign OE_DATA_52_const_net_2              = 4'h0;
assign OE_DATA_53_const_net_2              = 4'h0;
assign OE_DATA_54_const_net_2              = 4'h0;
assign OE_DATA_55_const_net_2              = 4'h0;
assign OE_DATA_56_const_net_2              = 4'h0;
assign OE_DATA_57_const_net_2              = 4'h0;
assign OE_DATA_58_const_net_2              = 4'h0;
assign OE_DATA_59_const_net_2              = 4'h0;
assign OE_DATA_60_const_net_2              = 4'h0;
assign OE_DATA_61_const_net_2              = 4'h0;
assign OE_DATA_62_const_net_2              = 4'h0;
assign OE_DATA_63_const_net_2              = 4'h0;
assign OE_DATA_64_const_net_2              = 4'h0;
assign OE_DATA_65_const_net_2              = 4'h0;
assign OE_DATA_66_const_net_2              = 4'h0;
assign OE_DATA_67_const_net_2              = 4'h0;
assign OE_DATA_68_const_net_2              = 4'h0;
assign OE_DATA_69_const_net_2              = 4'h0;
assign OE_DATA_70_const_net_2              = 4'h0;
assign OE_DATA_71_const_net_2              = 4'h0;
assign OE_DATA_72_const_net_2              = 4'h0;
assign OE_DATA_73_const_net_2              = 4'h0;
assign OE_DATA_74_const_net_2              = 4'h0;
assign OE_DATA_75_const_net_2              = 4'h0;
assign OE_DATA_76_const_net_2              = 4'h0;
assign OE_DATA_77_const_net_2              = 4'h0;
assign OE_DATA_78_const_net_2              = 4'h0;
assign OE_DATA_79_const_net_2              = 4'h0;
assign OE_DATA_80_const_net_2              = 4'h0;
assign OE_DATA_81_const_net_2              = 4'h0;
assign OE_DATA_82_const_net_2              = 4'h0;
assign OE_DATA_83_const_net_2              = 4'h0;
assign OE_DATA_84_const_net_2              = 4'h0;
assign OE_DATA_85_const_net_2              = 4'h0;
assign OE_DATA_86_const_net_2              = 4'h0;
assign OE_DATA_87_const_net_2              = 4'h0;
assign OE_DATA_88_const_net_2              = 4'h0;
assign OE_DATA_89_const_net_2              = 4'h0;
assign OE_DATA_90_const_net_2              = 4'h0;
assign OE_DATA_91_const_net_2              = 4'h0;
assign OE_DATA_92_const_net_2              = 4'h0;
assign OE_DATA_93_const_net_2              = 4'h0;
assign OE_DATA_94_const_net_2              = 4'h0;
assign OE_DATA_95_const_net_2              = 4'h0;
assign OE_DATA_96_const_net_2              = 4'h0;
assign OE_DATA_97_const_net_2              = 4'h0;
assign OE_DATA_98_const_net_2              = 4'h0;
assign OE_DATA_99_const_net_2              = 4'h0;
assign OE_DATA_100_const_net_2             = 4'h0;
assign OE_DATA_101_const_net_2             = 4'h0;
assign OE_DATA_102_const_net_2             = 4'h0;
assign OE_DATA_103_const_net_2             = 4'h0;
assign OE_DATA_104_const_net_2             = 4'h0;
assign OE_DATA_105_const_net_2             = 4'h0;
assign OE_DATA_106_const_net_2             = 4'h0;
assign OE_DATA_107_const_net_2             = 4'h0;
assign OE_DATA_108_const_net_2             = 4'h0;
assign OE_DATA_109_const_net_2             = 4'h0;
assign OE_DATA_110_const_net_2             = 4'h0;
assign OE_DATA_111_const_net_2             = 4'h0;
assign OE_DATA_112_const_net_2             = 4'h0;
assign OE_DATA_113_const_net_2             = 4'h0;
assign OE_DATA_114_const_net_2             = 4'h0;
assign OE_DATA_115_const_net_2             = 4'h0;
assign OE_DATA_116_const_net_2             = 4'h0;
assign OE_DATA_117_const_net_2             = 4'h0;
assign OE_DATA_118_const_net_2             = 4'h0;
assign OE_DATA_119_const_net_2             = 4'h0;
assign OE_DATA_120_const_net_2             = 4'h0;
assign OE_DATA_121_const_net_2             = 4'h0;
assign OE_DATA_122_const_net_2             = 4'h0;
assign OE_DATA_123_const_net_2             = 4'h0;
assign OE_DATA_124_const_net_2             = 4'h0;
assign OE_DATA_125_const_net_2             = 4'h0;
assign OE_DATA_126_const_net_2             = 4'h0;
assign OE_DATA_127_const_net_2             = 4'h0;
assign RX_DQS_90_const_net_3               = 2'h0;
assign FIFO_WR_PTR_const_net_3             = 3'h0;
assign FIFO_RD_PTR_const_net_3             = 3'h0;
assign EYE_MONITOR_LANE_WIDTH_const_net_3  = 3'h0;
assign TX_DATA_1_const_net_2               = 4'h0;
assign TX_DATA_2_const_net_2               = 4'h0;
assign TX_DATA_3_const_net_2               = 4'h0;
assign TX_DATA_4_const_net_2               = 4'h0;
assign TX_DATA_5_const_net_2               = 4'h0;
assign TX_DATA_6_const_net_2               = 4'h0;
assign TX_DATA_7_const_net_2               = 4'h0;
assign TX_DATA_8_const_net_2               = 4'h0;
assign TX_DATA_9_const_net_2               = 4'h0;
assign TX_DATA_10_const_net_2              = 4'h0;
assign TX_DATA_11_const_net_2              = 4'h0;
assign TX_DATA_12_const_net_3              = 4'h0;
assign TX_DATA_13_const_net_3              = 4'h0;
assign TX_DATA_14_const_net_3              = 4'h0;
assign TX_DATA_15_const_net_3              = 4'h0;
assign TX_DATA_16_const_net_3              = 4'h0;
assign TX_DATA_17_const_net_3              = 4'h0;
assign TX_DATA_18_const_net_3              = 4'h0;
assign TX_DATA_19_const_net_3              = 4'h0;
assign TX_DATA_20_const_net_3              = 4'h0;
assign TX_DATA_21_const_net_3              = 4'h0;
assign TX_DATA_22_const_net_3              = 4'h0;
assign TX_DATA_23_const_net_3              = 4'h0;
assign TX_DATA_24_const_net_3              = 4'h0;
assign TX_DATA_25_const_net_3              = 4'h0;
assign TX_DATA_26_const_net_3              = 4'h0;
assign TX_DATA_27_const_net_3              = 4'h0;
assign TX_DATA_28_const_net_3              = 4'h0;
assign TX_DATA_29_const_net_3              = 4'h0;
assign TX_DATA_30_const_net_3              = 4'h0;
assign TX_DATA_31_const_net_3              = 4'h0;
assign TX_DATA_32_const_net_3              = 4'h0;
assign TX_DATA_33_const_net_3              = 4'h0;
assign TX_DATA_34_const_net_3              = 4'h0;
assign TX_DATA_35_const_net_3              = 4'h0;
assign TX_DATA_36_const_net_3              = 4'h0;
assign TX_DATA_37_const_net_3              = 4'h0;
assign TX_DATA_38_const_net_3              = 4'h0;
assign TX_DATA_39_const_net_3              = 4'h0;
assign TX_DATA_40_const_net_3              = 4'h0;
assign TX_DATA_41_const_net_3              = 4'h0;
assign TX_DATA_42_const_net_3              = 4'h0;
assign TX_DATA_43_const_net_3              = 4'h0;
assign TX_DATA_44_const_net_3              = 4'h0;
assign TX_DATA_45_const_net_3              = 4'h0;
assign TX_DATA_46_const_net_3              = 4'h0;
assign TX_DATA_47_const_net_3              = 4'h0;
assign TX_DATA_48_const_net_3              = 4'h0;
assign TX_DATA_49_const_net_3              = 4'h0;
assign TX_DATA_50_const_net_3              = 4'h0;
assign TX_DATA_51_const_net_3              = 4'h0;
assign TX_DATA_52_const_net_3              = 4'h0;
assign TX_DATA_53_const_net_3              = 4'h0;
assign TX_DATA_54_const_net_3              = 4'h0;
assign TX_DATA_55_const_net_3              = 4'h0;
assign TX_DATA_56_const_net_3              = 4'h0;
assign TX_DATA_57_const_net_3              = 4'h0;
assign TX_DATA_58_const_net_3              = 4'h0;
assign TX_DATA_59_const_net_3              = 4'h0;
assign TX_DATA_60_const_net_3              = 4'h0;
assign TX_DATA_61_const_net_3              = 4'h0;
assign TX_DATA_62_const_net_3              = 4'h0;
assign TX_DATA_63_const_net_3              = 4'h0;
assign TX_DATA_64_const_net_3              = 4'h0;
assign TX_DATA_65_const_net_3              = 4'h0;
assign TX_DATA_66_const_net_3              = 4'h0;
assign TX_DATA_67_const_net_3              = 4'h0;
assign TX_DATA_68_const_net_3              = 4'h0;
assign TX_DATA_69_const_net_3              = 4'h0;
assign TX_DATA_70_const_net_3              = 4'h0;
assign TX_DATA_71_const_net_3              = 4'h0;
assign TX_DATA_72_const_net_3              = 4'h0;
assign TX_DATA_73_const_net_3              = 4'h0;
assign TX_DATA_74_const_net_3              = 4'h0;
assign TX_DATA_75_const_net_3              = 4'h0;
assign TX_DATA_76_const_net_3              = 4'h0;
assign TX_DATA_77_const_net_3              = 4'h0;
assign TX_DATA_78_const_net_3              = 4'h0;
assign TX_DATA_79_const_net_3              = 4'h0;
assign TX_DATA_80_const_net_3              = 4'h0;
assign TX_DATA_81_const_net_3              = 4'h0;
assign TX_DATA_82_const_net_3              = 4'h0;
assign TX_DATA_83_const_net_3              = 4'h0;
assign TX_DATA_84_const_net_3              = 4'h0;
assign TX_DATA_85_const_net_3              = 4'h0;
assign TX_DATA_86_const_net_3              = 4'h0;
assign TX_DATA_87_const_net_3              = 4'h0;
assign TX_DATA_88_const_net_3              = 4'h0;
assign TX_DATA_89_const_net_3              = 4'h0;
assign TX_DATA_90_const_net_3              = 4'h0;
assign TX_DATA_91_const_net_3              = 4'h0;
assign TX_DATA_92_const_net_3              = 4'h0;
assign TX_DATA_93_const_net_3              = 4'h0;
assign TX_DATA_94_const_net_3              = 4'h0;
assign TX_DATA_95_const_net_3              = 4'h0;
assign TX_DATA_96_const_net_3              = 4'h0;
assign TX_DATA_97_const_net_3              = 4'h0;
assign TX_DATA_98_const_net_3              = 4'h0;
assign TX_DATA_99_const_net_3              = 4'h0;
assign TX_DATA_100_const_net_3             = 4'h0;
assign TX_DATA_101_const_net_3             = 4'h0;
assign TX_DATA_102_const_net_3             = 4'h0;
assign TX_DATA_103_const_net_3             = 4'h0;
assign TX_DATA_104_const_net_3             = 4'h0;
assign TX_DATA_105_const_net_3             = 4'h0;
assign TX_DATA_106_const_net_3             = 4'h0;
assign TX_DATA_107_const_net_3             = 4'h0;
assign TX_DATA_108_const_net_3             = 4'h0;
assign TX_DATA_109_const_net_3             = 4'h0;
assign TX_DATA_110_const_net_3             = 4'h0;
assign TX_DATA_111_const_net_3             = 4'h0;
assign TX_DATA_112_const_net_3             = 4'h0;
assign TX_DATA_113_const_net_3             = 4'h0;
assign TX_DATA_114_const_net_3             = 4'h0;
assign TX_DATA_115_const_net_3             = 4'h0;
assign TX_DATA_116_const_net_3             = 4'h0;
assign TX_DATA_117_const_net_3             = 4'h0;
assign TX_DATA_118_const_net_3             = 4'h0;
assign TX_DATA_119_const_net_3             = 4'h0;
assign TX_DATA_120_const_net_3             = 4'h0;
assign TX_DATA_121_const_net_3             = 4'h0;
assign TX_DATA_122_const_net_3             = 4'h0;
assign TX_DATA_123_const_net_3             = 4'h0;
assign TX_DATA_124_const_net_3             = 4'h0;
assign TX_DATA_125_const_net_3             = 4'h0;
assign TX_DATA_126_const_net_3             = 4'h0;
assign TX_DATA_127_const_net_3             = 4'h0;
assign OE_DATA_1_const_net_5               = 4'h0;
assign OE_DATA_2_const_net_3               = 4'h0;
assign OE_DATA_3_const_net_3               = 4'h0;
assign OE_DATA_4_const_net_3               = 4'h0;
assign OE_DATA_5_const_net_3               = 4'h0;
assign OE_DATA_6_const_net_3               = 4'h0;
assign OE_DATA_7_const_net_3               = 4'h0;
assign OE_DATA_8_const_net_3               = 4'h0;
assign OE_DATA_9_const_net_3               = 4'h0;
assign OE_DATA_10_const_net_3              = 4'h0;
assign OE_DATA_11_const_net_3              = 4'h0;
assign OE_DATA_12_const_net_3              = 4'h0;
assign OE_DATA_13_const_net_3              = 4'h0;
assign OE_DATA_14_const_net_3              = 4'h0;
assign OE_DATA_15_const_net_3              = 4'h0;
assign OE_DATA_16_const_net_3              = 4'h0;
assign OE_DATA_17_const_net_3              = 4'h0;
assign OE_DATA_18_const_net_3              = 4'h0;
assign OE_DATA_19_const_net_3              = 4'h0;
assign OE_DATA_20_const_net_3              = 4'h0;
assign OE_DATA_21_const_net_3              = 4'h0;
assign OE_DATA_22_const_net_3              = 4'h0;
assign OE_DATA_23_const_net_3              = 4'h0;
assign OE_DATA_24_const_net_3              = 4'h0;
assign OE_DATA_25_const_net_3              = 4'h0;
assign OE_DATA_26_const_net_3              = 4'h0;
assign OE_DATA_27_const_net_3              = 4'h0;
assign OE_DATA_28_const_net_3              = 4'h0;
assign OE_DATA_29_const_net_3              = 4'h0;
assign OE_DATA_30_const_net_3              = 4'h0;
assign OE_DATA_31_const_net_3              = 4'h0;
assign OE_DATA_32_const_net_3              = 4'h0;
assign OE_DATA_33_const_net_3              = 4'h0;
assign OE_DATA_34_const_net_3              = 4'h0;
assign OE_DATA_35_const_net_3              = 4'h0;
assign OE_DATA_36_const_net_3              = 4'h0;
assign OE_DATA_37_const_net_3              = 4'h0;
assign OE_DATA_38_const_net_3              = 4'h0;
assign OE_DATA_39_const_net_3              = 4'h0;
assign OE_DATA_40_const_net_3              = 4'h0;
assign OE_DATA_41_const_net_3              = 4'h0;
assign OE_DATA_42_const_net_3              = 4'h0;
assign OE_DATA_43_const_net_3              = 4'h0;
assign OE_DATA_44_const_net_3              = 4'h0;
assign OE_DATA_45_const_net_3              = 4'h0;
assign OE_DATA_46_const_net_3              = 4'h0;
assign OE_DATA_47_const_net_3              = 4'h0;
assign OE_DATA_48_const_net_3              = 4'h0;
assign OE_DATA_49_const_net_3              = 4'h0;
assign OE_DATA_50_const_net_3              = 4'h0;
assign OE_DATA_51_const_net_3              = 4'h0;
assign OE_DATA_52_const_net_3              = 4'h0;
assign OE_DATA_53_const_net_3              = 4'h0;
assign OE_DATA_54_const_net_3              = 4'h0;
assign OE_DATA_55_const_net_3              = 4'h0;
assign OE_DATA_56_const_net_3              = 4'h0;
assign OE_DATA_57_const_net_3              = 4'h0;
assign OE_DATA_58_const_net_3              = 4'h0;
assign OE_DATA_59_const_net_3              = 4'h0;
assign OE_DATA_60_const_net_3              = 4'h0;
assign OE_DATA_61_const_net_3              = 4'h0;
assign OE_DATA_62_const_net_3              = 4'h0;
assign OE_DATA_63_const_net_3              = 4'h0;
assign OE_DATA_64_const_net_3              = 4'h0;
assign OE_DATA_65_const_net_3              = 4'h0;
assign OE_DATA_66_const_net_3              = 4'h0;
assign OE_DATA_67_const_net_3              = 4'h0;
assign OE_DATA_68_const_net_3              = 4'h0;
assign OE_DATA_69_const_net_3              = 4'h0;
assign OE_DATA_70_const_net_3              = 4'h0;
assign OE_DATA_71_const_net_3              = 4'h0;
assign OE_DATA_72_const_net_3              = 4'h0;
assign OE_DATA_73_const_net_3              = 4'h0;
assign OE_DATA_74_const_net_3              = 4'h0;
assign OE_DATA_75_const_net_3              = 4'h0;
assign OE_DATA_76_const_net_3              = 4'h0;
assign OE_DATA_77_const_net_3              = 4'h0;
assign OE_DATA_78_const_net_3              = 4'h0;
assign OE_DATA_79_const_net_3              = 4'h0;
assign OE_DATA_80_const_net_3              = 4'h0;
assign OE_DATA_81_const_net_3              = 4'h0;
assign OE_DATA_82_const_net_3              = 4'h0;
assign OE_DATA_83_const_net_3              = 4'h0;
assign OE_DATA_84_const_net_3              = 4'h0;
assign OE_DATA_85_const_net_3              = 4'h0;
assign OE_DATA_86_const_net_3              = 4'h0;
assign OE_DATA_87_const_net_3              = 4'h0;
assign OE_DATA_88_const_net_3              = 4'h0;
assign OE_DATA_89_const_net_3              = 4'h0;
assign OE_DATA_90_const_net_3              = 4'h0;
assign OE_DATA_91_const_net_3              = 4'h0;
assign OE_DATA_92_const_net_3              = 4'h0;
assign OE_DATA_93_const_net_3              = 4'h0;
assign OE_DATA_94_const_net_3              = 4'h0;
assign OE_DATA_95_const_net_3              = 4'h0;
assign OE_DATA_96_const_net_3              = 4'h0;
assign OE_DATA_97_const_net_3              = 4'h0;
assign OE_DATA_98_const_net_3              = 4'h0;
assign OE_DATA_99_const_net_3              = 4'h0;
assign OE_DATA_100_const_net_3             = 4'h0;
assign OE_DATA_101_const_net_3             = 4'h0;
assign OE_DATA_102_const_net_3             = 4'h0;
assign OE_DATA_103_const_net_3             = 4'h0;
assign OE_DATA_104_const_net_3             = 4'h0;
assign OE_DATA_105_const_net_3             = 4'h0;
assign OE_DATA_106_const_net_3             = 4'h0;
assign OE_DATA_107_const_net_3             = 4'h0;
assign OE_DATA_108_const_net_3             = 4'h0;
assign OE_DATA_109_const_net_3             = 4'h0;
assign OE_DATA_110_const_net_3             = 4'h0;
assign OE_DATA_111_const_net_3             = 4'h0;
assign OE_DATA_112_const_net_3             = 4'h0;
assign OE_DATA_113_const_net_3             = 4'h0;
assign OE_DATA_114_const_net_3             = 4'h0;
assign OE_DATA_115_const_net_3             = 4'h0;
assign OE_DATA_116_const_net_3             = 4'h0;
assign OE_DATA_117_const_net_3             = 4'h0;
assign OE_DATA_118_const_net_3             = 4'h0;
assign OE_DATA_119_const_net_3             = 4'h0;
assign OE_DATA_120_const_net_3             = 4'h0;
assign OE_DATA_121_const_net_3             = 4'h0;
assign OE_DATA_122_const_net_3             = 4'h0;
assign OE_DATA_123_const_net_3             = 4'h0;
assign OE_DATA_124_const_net_3             = 4'h0;
assign OE_DATA_125_const_net_3             = 4'h0;
assign OE_DATA_126_const_net_3             = 4'h0;
assign OE_DATA_127_const_net_3             = 4'h0;
assign RX_DQS_90_const_net_4               = 2'h0;
assign FIFO_WR_PTR_const_net_4             = 3'h0;
assign FIFO_RD_PTR_const_net_4             = 3'h0;
assign EYE_MONITOR_LANE_WIDTH_const_net_4  = 3'h0;
assign TX_DATA_2_const_net_3               = 4'h0;
assign TX_DATA_3_const_net_3               = 4'h0;
assign TX_DATA_4_const_net_3               = 4'h0;
assign TX_DATA_5_const_net_3               = 4'h0;
assign TX_DATA_6_const_net_3               = 4'h0;
assign TX_DATA_7_const_net_3               = 4'h0;
assign TX_DATA_8_const_net_3               = 4'h0;
assign TX_DATA_9_const_net_3               = 4'h0;
assign TX_DATA_10_const_net_3              = 4'h0;
assign TX_DATA_11_const_net_3              = 4'h0;
assign TX_DATA_12_const_net_4              = 4'h0;
assign TX_DATA_13_const_net_4              = 4'h0;
assign TX_DATA_14_const_net_4              = 4'h0;
assign TX_DATA_15_const_net_4              = 4'h0;
assign TX_DATA_16_const_net_4              = 4'h0;
assign TX_DATA_17_const_net_4              = 4'h0;
assign TX_DATA_18_const_net_4              = 4'h0;
assign TX_DATA_19_const_net_4              = 4'h0;
assign TX_DATA_20_const_net_4              = 4'h0;
assign TX_DATA_21_const_net_4              = 4'h0;
assign TX_DATA_22_const_net_4              = 4'h0;
assign TX_DATA_23_const_net_4              = 4'h0;
assign TX_DATA_24_const_net_4              = 4'h0;
assign TX_DATA_25_const_net_4              = 4'h0;
assign TX_DATA_26_const_net_4              = 4'h0;
assign TX_DATA_27_const_net_4              = 4'h0;
assign TX_DATA_28_const_net_4              = 4'h0;
assign TX_DATA_29_const_net_4              = 4'h0;
assign TX_DATA_30_const_net_4              = 4'h0;
assign TX_DATA_31_const_net_4              = 4'h0;
assign TX_DATA_32_const_net_4              = 4'h0;
assign TX_DATA_33_const_net_4              = 4'h0;
assign TX_DATA_34_const_net_4              = 4'h0;
assign TX_DATA_35_const_net_4              = 4'h0;
assign TX_DATA_36_const_net_4              = 4'h0;
assign TX_DATA_37_const_net_4              = 4'h0;
assign TX_DATA_38_const_net_4              = 4'h0;
assign TX_DATA_39_const_net_4              = 4'h0;
assign TX_DATA_40_const_net_4              = 4'h0;
assign TX_DATA_41_const_net_4              = 4'h0;
assign TX_DATA_42_const_net_4              = 4'h0;
assign TX_DATA_43_const_net_4              = 4'h0;
assign TX_DATA_44_const_net_4              = 4'h0;
assign TX_DATA_45_const_net_4              = 4'h0;
assign TX_DATA_46_const_net_4              = 4'h0;
assign TX_DATA_47_const_net_4              = 4'h0;
assign TX_DATA_48_const_net_4              = 4'h0;
assign TX_DATA_49_const_net_4              = 4'h0;
assign TX_DATA_50_const_net_4              = 4'h0;
assign TX_DATA_51_const_net_4              = 4'h0;
assign TX_DATA_52_const_net_4              = 4'h0;
assign TX_DATA_53_const_net_4              = 4'h0;
assign TX_DATA_54_const_net_4              = 4'h0;
assign TX_DATA_55_const_net_4              = 4'h0;
assign TX_DATA_56_const_net_4              = 4'h0;
assign TX_DATA_57_const_net_4              = 4'h0;
assign TX_DATA_58_const_net_4              = 4'h0;
assign TX_DATA_59_const_net_4              = 4'h0;
assign TX_DATA_60_const_net_4              = 4'h0;
assign TX_DATA_61_const_net_4              = 4'h0;
assign TX_DATA_62_const_net_4              = 4'h0;
assign TX_DATA_63_const_net_4              = 4'h0;
assign TX_DATA_64_const_net_4              = 4'h0;
assign TX_DATA_65_const_net_4              = 4'h0;
assign TX_DATA_66_const_net_4              = 4'h0;
assign TX_DATA_67_const_net_4              = 4'h0;
assign TX_DATA_68_const_net_4              = 4'h0;
assign TX_DATA_69_const_net_4              = 4'h0;
assign TX_DATA_70_const_net_4              = 4'h0;
assign TX_DATA_71_const_net_4              = 4'h0;
assign TX_DATA_72_const_net_4              = 4'h0;
assign TX_DATA_73_const_net_4              = 4'h0;
assign TX_DATA_74_const_net_4              = 4'h0;
assign TX_DATA_75_const_net_4              = 4'h0;
assign TX_DATA_76_const_net_4              = 4'h0;
assign TX_DATA_77_const_net_4              = 4'h0;
assign TX_DATA_78_const_net_4              = 4'h0;
assign TX_DATA_79_const_net_4              = 4'h0;
assign TX_DATA_80_const_net_4              = 4'h0;
assign TX_DATA_81_const_net_4              = 4'h0;
assign TX_DATA_82_const_net_4              = 4'h0;
assign TX_DATA_83_const_net_4              = 4'h0;
assign TX_DATA_84_const_net_4              = 4'h0;
assign TX_DATA_85_const_net_4              = 4'h0;
assign TX_DATA_86_const_net_4              = 4'h0;
assign TX_DATA_87_const_net_4              = 4'h0;
assign TX_DATA_88_const_net_4              = 4'h0;
assign TX_DATA_89_const_net_4              = 4'h0;
assign TX_DATA_90_const_net_4              = 4'h0;
assign TX_DATA_91_const_net_4              = 4'h0;
assign TX_DATA_92_const_net_4              = 4'h0;
assign TX_DATA_93_const_net_4              = 4'h0;
assign TX_DATA_94_const_net_4              = 4'h0;
assign TX_DATA_95_const_net_4              = 4'h0;
assign TX_DATA_96_const_net_4              = 4'h0;
assign TX_DATA_97_const_net_4              = 4'h0;
assign TX_DATA_98_const_net_4              = 4'h0;
assign TX_DATA_99_const_net_4              = 4'h0;
assign TX_DATA_100_const_net_4             = 4'h0;
assign TX_DATA_101_const_net_4             = 4'h0;
assign TX_DATA_102_const_net_4             = 4'h0;
assign TX_DATA_103_const_net_4             = 4'h0;
assign TX_DATA_104_const_net_4             = 4'h0;
assign TX_DATA_105_const_net_4             = 4'h0;
assign TX_DATA_106_const_net_4             = 4'h0;
assign TX_DATA_107_const_net_4             = 4'h0;
assign TX_DATA_108_const_net_4             = 4'h0;
assign TX_DATA_109_const_net_4             = 4'h0;
assign TX_DATA_110_const_net_4             = 4'h0;
assign TX_DATA_111_const_net_4             = 4'h0;
assign TX_DATA_112_const_net_4             = 4'h0;
assign TX_DATA_113_const_net_4             = 4'h0;
assign TX_DATA_114_const_net_4             = 4'h0;
assign TX_DATA_115_const_net_4             = 4'h0;
assign TX_DATA_116_const_net_4             = 4'h0;
assign TX_DATA_117_const_net_4             = 4'h0;
assign TX_DATA_118_const_net_4             = 4'h0;
assign TX_DATA_119_const_net_4             = 4'h0;
assign TX_DATA_120_const_net_4             = 4'h0;
assign TX_DATA_121_const_net_4             = 4'h0;
assign TX_DATA_122_const_net_4             = 4'h0;
assign TX_DATA_123_const_net_4             = 4'h0;
assign TX_DATA_124_const_net_4             = 4'h0;
assign TX_DATA_125_const_net_4             = 4'h0;
assign TX_DATA_126_const_net_4             = 4'h0;
assign TX_DATA_127_const_net_4             = 4'h0;
assign OE_DATA_2_const_net_4               = 4'h0;
assign OE_DATA_3_const_net_4               = 4'h0;
assign OE_DATA_4_const_net_4               = 4'h0;
assign OE_DATA_5_const_net_4               = 4'h0;
assign OE_DATA_6_const_net_4               = 4'h0;
assign OE_DATA_7_const_net_4               = 4'h0;
assign OE_DATA_8_const_net_4               = 4'h0;
assign OE_DATA_9_const_net_4               = 4'h0;
assign OE_DATA_10_const_net_4              = 4'h0;
assign OE_DATA_11_const_net_4              = 4'h0;
assign OE_DATA_12_const_net_4              = 4'h0;
assign OE_DATA_13_const_net_4              = 4'h0;
assign OE_DATA_14_const_net_4              = 4'h0;
assign OE_DATA_15_const_net_4              = 4'h0;
assign OE_DATA_16_const_net_4              = 4'h0;
assign OE_DATA_17_const_net_4              = 4'h0;
assign OE_DATA_18_const_net_4              = 4'h0;
assign OE_DATA_19_const_net_4              = 4'h0;
assign OE_DATA_20_const_net_4              = 4'h0;
assign OE_DATA_21_const_net_4              = 4'h0;
assign OE_DATA_22_const_net_4              = 4'h0;
assign OE_DATA_23_const_net_4              = 4'h0;
assign OE_DATA_24_const_net_4              = 4'h0;
assign OE_DATA_25_const_net_4              = 4'h0;
assign OE_DATA_26_const_net_4              = 4'h0;
assign OE_DATA_27_const_net_4              = 4'h0;
assign OE_DATA_28_const_net_4              = 4'h0;
assign OE_DATA_29_const_net_4              = 4'h0;
assign OE_DATA_30_const_net_4              = 4'h0;
assign OE_DATA_31_const_net_4              = 4'h0;
assign OE_DATA_32_const_net_4              = 4'h0;
assign OE_DATA_33_const_net_4              = 4'h0;
assign OE_DATA_34_const_net_4              = 4'h0;
assign OE_DATA_35_const_net_4              = 4'h0;
assign OE_DATA_36_const_net_4              = 4'h0;
assign OE_DATA_37_const_net_4              = 4'h0;
assign OE_DATA_38_const_net_4              = 4'h0;
assign OE_DATA_39_const_net_4              = 4'h0;
assign OE_DATA_40_const_net_4              = 4'h0;
assign OE_DATA_41_const_net_4              = 4'h0;
assign OE_DATA_42_const_net_4              = 4'h0;
assign OE_DATA_43_const_net_4              = 4'h0;
assign OE_DATA_44_const_net_4              = 4'h0;
assign OE_DATA_45_const_net_4              = 4'h0;
assign OE_DATA_46_const_net_4              = 4'h0;
assign OE_DATA_47_const_net_4              = 4'h0;
assign OE_DATA_48_const_net_4              = 4'h0;
assign OE_DATA_49_const_net_4              = 4'h0;
assign OE_DATA_50_const_net_4              = 4'h0;
assign OE_DATA_51_const_net_4              = 4'h0;
assign OE_DATA_52_const_net_4              = 4'h0;
assign OE_DATA_53_const_net_4              = 4'h0;
assign OE_DATA_54_const_net_4              = 4'h0;
assign OE_DATA_55_const_net_4              = 4'h0;
assign OE_DATA_56_const_net_4              = 4'h0;
assign OE_DATA_57_const_net_4              = 4'h0;
assign OE_DATA_58_const_net_4              = 4'h0;
assign OE_DATA_59_const_net_4              = 4'h0;
assign OE_DATA_60_const_net_4              = 4'h0;
assign OE_DATA_61_const_net_4              = 4'h0;
assign OE_DATA_62_const_net_4              = 4'h0;
assign OE_DATA_63_const_net_4              = 4'h0;
assign OE_DATA_64_const_net_4              = 4'h0;
assign OE_DATA_65_const_net_4              = 4'h0;
assign OE_DATA_66_const_net_4              = 4'h0;
assign OE_DATA_67_const_net_4              = 4'h0;
assign OE_DATA_68_const_net_4              = 4'h0;
assign OE_DATA_69_const_net_4              = 4'h0;
assign OE_DATA_70_const_net_4              = 4'h0;
assign OE_DATA_71_const_net_4              = 4'h0;
assign OE_DATA_72_const_net_4              = 4'h0;
assign OE_DATA_73_const_net_4              = 4'h0;
assign OE_DATA_74_const_net_4              = 4'h0;
assign OE_DATA_75_const_net_4              = 4'h0;
assign OE_DATA_76_const_net_4              = 4'h0;
assign OE_DATA_77_const_net_4              = 4'h0;
assign OE_DATA_78_const_net_4              = 4'h0;
assign OE_DATA_79_const_net_4              = 4'h0;
assign OE_DATA_80_const_net_4              = 4'h0;
assign OE_DATA_81_const_net_4              = 4'h0;
assign OE_DATA_82_const_net_4              = 4'h0;
assign OE_DATA_83_const_net_4              = 4'h0;
assign OE_DATA_84_const_net_4              = 4'h0;
assign OE_DATA_85_const_net_4              = 4'h0;
assign OE_DATA_86_const_net_4              = 4'h0;
assign OE_DATA_87_const_net_4              = 4'h0;
assign OE_DATA_88_const_net_4              = 4'h0;
assign OE_DATA_89_const_net_4              = 4'h0;
assign OE_DATA_90_const_net_4              = 4'h0;
assign OE_DATA_91_const_net_4              = 4'h0;
assign OE_DATA_92_const_net_4              = 4'h0;
assign OE_DATA_93_const_net_4              = 4'h0;
assign OE_DATA_94_const_net_4              = 4'h0;
assign OE_DATA_95_const_net_4              = 4'h0;
assign OE_DATA_96_const_net_4              = 4'h0;
assign OE_DATA_97_const_net_4              = 4'h0;
assign OE_DATA_98_const_net_4              = 4'h0;
assign OE_DATA_99_const_net_4              = 4'h0;
assign OE_DATA_100_const_net_4             = 4'h0;
assign OE_DATA_101_const_net_4             = 4'h0;
assign OE_DATA_102_const_net_4             = 4'h0;
assign OE_DATA_103_const_net_4             = 4'h0;
assign OE_DATA_104_const_net_4             = 4'h0;
assign OE_DATA_105_const_net_4             = 4'h0;
assign OE_DATA_106_const_net_4             = 4'h0;
assign OE_DATA_107_const_net_4             = 4'h0;
assign OE_DATA_108_const_net_4             = 4'h0;
assign OE_DATA_109_const_net_4             = 4'h0;
assign OE_DATA_110_const_net_4             = 4'h0;
assign OE_DATA_111_const_net_4             = 4'h0;
assign OE_DATA_112_const_net_4             = 4'h0;
assign OE_DATA_113_const_net_4             = 4'h0;
assign OE_DATA_114_const_net_4             = 4'h0;
assign OE_DATA_115_const_net_4             = 4'h0;
assign OE_DATA_116_const_net_4             = 4'h0;
assign OE_DATA_117_const_net_4             = 4'h0;
assign OE_DATA_118_const_net_4             = 4'h0;
assign OE_DATA_119_const_net_4             = 4'h0;
assign OE_DATA_120_const_net_4             = 4'h0;
assign OE_DATA_121_const_net_4             = 4'h0;
assign OE_DATA_122_const_net_4             = 4'h0;
assign OE_DATA_123_const_net_4             = 4'h0;
assign OE_DATA_124_const_net_4             = 4'h0;
assign OE_DATA_125_const_net_4             = 4'h0;
assign OE_DATA_126_const_net_4             = 4'h0;
assign OE_DATA_127_const_net_4             = 4'h0;
assign PAD_const_net_1                     = 2'h0;
assign PAD_I_const_net_1                   = 2'h0;
assign PAD_N_const_net_1                   = 2'h0;
assign PAD_I_N_const_net_1                 = 2'h0;
assign RX_DQS_90_const_net_5               = 2'h0;
assign FIFO_WR_PTR_const_net_5             = 3'h0;
assign FIFO_RD_PTR_const_net_5             = 3'h0;
assign EYE_MONITOR_LANE_WIDTH_const_net_5  = 3'h0;
assign TX_DATA_0_const_net_8               = 8'h00;
assign TX_DATA_1_const_net_3               = 8'h00;
assign TX_DATA_2_const_net_4               = 8'h00;
assign TX_DATA_3_const_net_4               = 8'h00;
assign TX_DATA_4_const_net_4               = 8'h00;
assign TX_DATA_5_const_net_4               = 8'h00;
assign TX_DATA_6_const_net_4               = 8'h00;
assign TX_DATA_7_const_net_4               = 8'h00;
assign TX_DATA_8_const_net_4               = 8'h00;
assign TX_DATA_9_const_net_4               = 8'h00;
assign TX_DATA_10_const_net_4              = 8'h00;
assign TX_DATA_11_const_net_4              = 8'h00;
assign TX_DATA_12_const_net_5              = 8'h00;
assign TX_DATA_13_const_net_5              = 8'h00;
assign TX_DATA_14_const_net_5              = 8'h00;
assign TX_DATA_15_const_net_5              = 8'h00;
assign TX_DATA_16_const_net_5              = 8'h00;
assign TX_DATA_17_const_net_5              = 8'h00;
assign TX_DATA_18_const_net_5              = 8'h00;
assign TX_DATA_19_const_net_5              = 8'h00;
assign TX_DATA_20_const_net_5              = 8'h00;
assign TX_DATA_21_const_net_5              = 8'h00;
assign TX_DATA_22_const_net_5              = 8'h00;
assign TX_DATA_23_const_net_5              = 8'h00;
assign TX_DATA_24_const_net_5              = 8'h00;
assign TX_DATA_25_const_net_5              = 8'h00;
assign TX_DATA_26_const_net_5              = 8'h00;
assign TX_DATA_27_const_net_5              = 8'h00;
assign TX_DATA_28_const_net_5              = 8'h00;
assign TX_DATA_29_const_net_5              = 8'h00;
assign TX_DATA_30_const_net_5              = 8'h00;
assign TX_DATA_31_const_net_5              = 8'h00;
assign TX_DATA_32_const_net_5              = 8'h00;
assign TX_DATA_33_const_net_5              = 8'h00;
assign TX_DATA_34_const_net_5              = 8'h00;
assign TX_DATA_35_const_net_5              = 8'h00;
assign TX_DATA_36_const_net_5              = 8'h00;
assign TX_DATA_37_const_net_5              = 8'h00;
assign TX_DATA_38_const_net_5              = 8'h00;
assign TX_DATA_39_const_net_5              = 8'h00;
assign TX_DATA_40_const_net_5              = 8'h00;
assign TX_DATA_41_const_net_5              = 8'h00;
assign TX_DATA_42_const_net_5              = 8'h00;
assign TX_DATA_43_const_net_5              = 8'h00;
assign TX_DATA_44_const_net_5              = 8'h00;
assign TX_DATA_45_const_net_5              = 8'h00;
assign TX_DATA_46_const_net_5              = 8'h00;
assign TX_DATA_47_const_net_5              = 8'h00;
assign TX_DATA_48_const_net_5              = 8'h00;
assign TX_DATA_49_const_net_5              = 8'h00;
assign TX_DATA_50_const_net_5              = 8'h00;
assign TX_DATA_51_const_net_5              = 8'h00;
assign TX_DATA_52_const_net_5              = 8'h00;
assign TX_DATA_53_const_net_5              = 8'h00;
assign TX_DATA_54_const_net_5              = 8'h00;
assign TX_DATA_55_const_net_5              = 8'h00;
assign TX_DATA_56_const_net_5              = 8'h00;
assign TX_DATA_57_const_net_5              = 8'h00;
assign TX_DATA_58_const_net_5              = 8'h00;
assign TX_DATA_59_const_net_5              = 8'h00;
assign TX_DATA_60_const_net_5              = 8'h00;
assign TX_DATA_61_const_net_5              = 8'h00;
assign TX_DATA_62_const_net_5              = 8'h00;
assign TX_DATA_63_const_net_5              = 8'h00;
assign TX_DATA_64_const_net_5              = 8'h00;
assign TX_DATA_65_const_net_5              = 8'h00;
assign TX_DATA_66_const_net_5              = 8'h00;
assign TX_DATA_67_const_net_5              = 8'h00;
assign TX_DATA_68_const_net_5              = 8'h00;
assign TX_DATA_69_const_net_5              = 8'h00;
assign TX_DATA_70_const_net_5              = 8'h00;
assign TX_DATA_71_const_net_5              = 8'h00;
assign TX_DATA_72_const_net_5              = 8'h00;
assign TX_DATA_73_const_net_5              = 8'h00;
assign TX_DATA_74_const_net_5              = 8'h00;
assign TX_DATA_75_const_net_5              = 8'h00;
assign TX_DATA_76_const_net_5              = 8'h00;
assign TX_DATA_77_const_net_5              = 8'h00;
assign TX_DATA_78_const_net_5              = 8'h00;
assign TX_DATA_79_const_net_5              = 8'h00;
assign TX_DATA_80_const_net_5              = 8'h00;
assign TX_DATA_81_const_net_5              = 8'h00;
assign TX_DATA_82_const_net_5              = 8'h00;
assign TX_DATA_83_const_net_5              = 8'h00;
assign TX_DATA_84_const_net_5              = 8'h00;
assign TX_DATA_85_const_net_5              = 8'h00;
assign TX_DATA_86_const_net_5              = 8'h00;
assign TX_DATA_87_const_net_5              = 8'h00;
assign TX_DATA_88_const_net_5              = 8'h00;
assign TX_DATA_89_const_net_5              = 8'h00;
assign TX_DATA_90_const_net_5              = 8'h00;
assign TX_DATA_91_const_net_5              = 8'h00;
assign TX_DATA_92_const_net_5              = 8'h00;
assign TX_DATA_93_const_net_5              = 8'h00;
assign TX_DATA_94_const_net_5              = 8'h00;
assign TX_DATA_95_const_net_5              = 8'h00;
assign TX_DATA_96_const_net_5              = 8'h00;
assign TX_DATA_97_const_net_5              = 8'h00;
assign TX_DATA_98_const_net_5              = 8'h00;
assign TX_DATA_99_const_net_5              = 8'h00;
assign TX_DATA_100_const_net_5             = 8'h00;
assign TX_DATA_101_const_net_5             = 8'h00;
assign TX_DATA_102_const_net_5             = 8'h00;
assign TX_DATA_103_const_net_5             = 8'h00;
assign TX_DATA_104_const_net_5             = 8'h00;
assign TX_DATA_105_const_net_5             = 8'h00;
assign TX_DATA_106_const_net_5             = 8'h00;
assign TX_DATA_107_const_net_5             = 8'h00;
assign TX_DATA_108_const_net_5             = 8'h00;
assign TX_DATA_109_const_net_5             = 8'h00;
assign TX_DATA_110_const_net_5             = 8'h00;
assign TX_DATA_111_const_net_5             = 8'h00;
assign TX_DATA_112_const_net_5             = 8'h00;
assign TX_DATA_113_const_net_5             = 8'h00;
assign TX_DATA_114_const_net_5             = 8'h00;
assign TX_DATA_115_const_net_5             = 8'h00;
assign TX_DATA_116_const_net_5             = 8'h00;
assign TX_DATA_117_const_net_5             = 8'h00;
assign TX_DATA_118_const_net_5             = 8'h00;
assign TX_DATA_119_const_net_5             = 8'h00;
assign TX_DATA_120_const_net_5             = 8'h00;
assign TX_DATA_121_const_net_5             = 8'h00;
assign TX_DATA_122_const_net_5             = 8'h00;
assign TX_DATA_123_const_net_5             = 8'h00;
assign TX_DATA_124_const_net_5             = 8'h00;
assign TX_DATA_125_const_net_5             = 8'h00;
assign TX_DATA_126_const_net_5             = 8'h00;
assign TX_DATA_127_const_net_5             = 8'h00;
assign OE_DATA_0_const_net_16              = 4'h0;
assign OE_DATA_1_const_net_6               = 4'h0;
assign OE_DATA_2_const_net_5               = 4'h0;
assign OE_DATA_3_const_net_5               = 4'h0;
assign OE_DATA_4_const_net_5               = 4'h0;
assign OE_DATA_5_const_net_5               = 4'h0;
assign OE_DATA_6_const_net_5               = 4'h0;
assign OE_DATA_7_const_net_5               = 4'h0;
assign OE_DATA_8_const_net_5               = 4'h0;
assign OE_DATA_9_const_net_5               = 4'h0;
assign OE_DATA_10_const_net_5              = 4'h0;
assign OE_DATA_11_const_net_5              = 4'h0;
assign OE_DATA_12_const_net_5              = 4'h0;
assign OE_DATA_13_const_net_5              = 4'h0;
assign OE_DATA_14_const_net_5              = 4'h0;
assign OE_DATA_15_const_net_5              = 4'h0;
assign OE_DATA_16_const_net_5              = 4'h0;
assign OE_DATA_17_const_net_5              = 4'h0;
assign OE_DATA_18_const_net_5              = 4'h0;
assign OE_DATA_19_const_net_5              = 4'h0;
assign OE_DATA_20_const_net_5              = 4'h0;
assign OE_DATA_21_const_net_5              = 4'h0;
assign OE_DATA_22_const_net_5              = 4'h0;
assign OE_DATA_23_const_net_5              = 4'h0;
assign OE_DATA_24_const_net_5              = 4'h0;
assign OE_DATA_25_const_net_5              = 4'h0;
assign OE_DATA_26_const_net_5              = 4'h0;
assign OE_DATA_27_const_net_5              = 4'h0;
assign OE_DATA_28_const_net_5              = 4'h0;
assign OE_DATA_29_const_net_5              = 4'h0;
assign OE_DATA_30_const_net_5              = 4'h0;
assign OE_DATA_31_const_net_5              = 4'h0;
assign OE_DATA_32_const_net_5              = 4'h0;
assign OE_DATA_33_const_net_5              = 4'h0;
assign OE_DATA_34_const_net_5              = 4'h0;
assign OE_DATA_35_const_net_5              = 4'h0;
assign OE_DATA_36_const_net_5              = 4'h0;
assign OE_DATA_37_const_net_5              = 4'h0;
assign OE_DATA_38_const_net_5              = 4'h0;
assign OE_DATA_39_const_net_5              = 4'h0;
assign OE_DATA_40_const_net_5              = 4'h0;
assign OE_DATA_41_const_net_5              = 4'h0;
assign OE_DATA_42_const_net_5              = 4'h0;
assign OE_DATA_43_const_net_5              = 4'h0;
assign OE_DATA_44_const_net_5              = 4'h0;
assign OE_DATA_45_const_net_5              = 4'h0;
assign OE_DATA_46_const_net_5              = 4'h0;
assign OE_DATA_47_const_net_5              = 4'h0;
assign OE_DATA_48_const_net_5              = 4'h0;
assign OE_DATA_49_const_net_5              = 4'h0;
assign OE_DATA_50_const_net_5              = 4'h0;
assign OE_DATA_51_const_net_5              = 4'h0;
assign OE_DATA_52_const_net_5              = 4'h0;
assign OE_DATA_53_const_net_5              = 4'h0;
assign OE_DATA_54_const_net_5              = 4'h0;
assign OE_DATA_55_const_net_5              = 4'h0;
assign OE_DATA_56_const_net_5              = 4'h0;
assign OE_DATA_57_const_net_5              = 4'h0;
assign OE_DATA_58_const_net_5              = 4'h0;
assign OE_DATA_59_const_net_5              = 4'h0;
assign OE_DATA_60_const_net_5              = 4'h0;
assign OE_DATA_61_const_net_5              = 4'h0;
assign OE_DATA_62_const_net_5              = 4'h0;
assign OE_DATA_63_const_net_5              = 4'h0;
assign OE_DATA_64_const_net_5              = 4'h0;
assign OE_DATA_65_const_net_5              = 4'h0;
assign OE_DATA_66_const_net_5              = 4'h0;
assign OE_DATA_67_const_net_5              = 4'h0;
assign OE_DATA_68_const_net_5              = 4'h0;
assign OE_DATA_69_const_net_5              = 4'h0;
assign OE_DATA_70_const_net_5              = 4'h0;
assign OE_DATA_71_const_net_5              = 4'h0;
assign OE_DATA_72_const_net_5              = 4'h0;
assign OE_DATA_73_const_net_5              = 4'h0;
assign OE_DATA_74_const_net_5              = 4'h0;
assign OE_DATA_75_const_net_5              = 4'h0;
assign OE_DATA_76_const_net_5              = 4'h0;
assign OE_DATA_77_const_net_5              = 4'h0;
assign OE_DATA_78_const_net_5              = 4'h0;
assign OE_DATA_79_const_net_5              = 4'h0;
assign OE_DATA_80_const_net_5              = 4'h0;
assign OE_DATA_81_const_net_5              = 4'h0;
assign OE_DATA_82_const_net_5              = 4'h0;
assign OE_DATA_83_const_net_5              = 4'h0;
assign OE_DATA_84_const_net_5              = 4'h0;
assign OE_DATA_85_const_net_5              = 4'h0;
assign OE_DATA_86_const_net_5              = 4'h0;
assign OE_DATA_87_const_net_5              = 4'h0;
assign OE_DATA_88_const_net_5              = 4'h0;
assign OE_DATA_89_const_net_5              = 4'h0;
assign OE_DATA_90_const_net_5              = 4'h0;
assign OE_DATA_91_const_net_5              = 4'h0;
assign OE_DATA_92_const_net_5              = 4'h0;
assign OE_DATA_93_const_net_5              = 4'h0;
assign OE_DATA_94_const_net_5              = 4'h0;
assign OE_DATA_95_const_net_5              = 4'h0;
assign OE_DATA_96_const_net_5              = 4'h0;
assign OE_DATA_97_const_net_5              = 4'h0;
assign OE_DATA_98_const_net_5              = 4'h0;
assign OE_DATA_99_const_net_5              = 4'h0;
assign OE_DATA_100_const_net_5             = 4'h0;
assign OE_DATA_101_const_net_5             = 4'h0;
assign OE_DATA_102_const_net_5             = 4'h0;
assign OE_DATA_103_const_net_5             = 4'h0;
assign OE_DATA_104_const_net_5             = 4'h0;
assign OE_DATA_105_const_net_5             = 4'h0;
assign OE_DATA_106_const_net_5             = 4'h0;
assign OE_DATA_107_const_net_5             = 4'h0;
assign OE_DATA_108_const_net_5             = 4'h0;
assign OE_DATA_109_const_net_5             = 4'h0;
assign OE_DATA_110_const_net_5             = 4'h0;
assign OE_DATA_111_const_net_5             = 4'h0;
assign OE_DATA_112_const_net_5             = 4'h0;
assign OE_DATA_113_const_net_5             = 4'h0;
assign OE_DATA_114_const_net_5             = 4'h0;
assign OE_DATA_115_const_net_5             = 4'h0;
assign OE_DATA_116_const_net_5             = 4'h0;
assign OE_DATA_117_const_net_5             = 4'h0;
assign OE_DATA_118_const_net_5             = 4'h0;
assign OE_DATA_119_const_net_5             = 4'h0;
assign OE_DATA_120_const_net_5             = 4'h0;
assign OE_DATA_121_const_net_5             = 4'h0;
assign OE_DATA_122_const_net_5             = 4'h0;
assign OE_DATA_123_const_net_5             = 4'h0;
assign OE_DATA_124_const_net_5             = 4'h0;
assign OE_DATA_125_const_net_5             = 4'h0;
assign OE_DATA_126_const_net_5             = 4'h0;
assign OE_DATA_127_const_net_5             = 4'h0;
assign RX_DQS_90_const_net_6               = 2'h0;
assign FIFO_WR_PTR_const_net_6             = 3'h0;
assign FIFO_RD_PTR_const_net_6             = 3'h0;
assign EYE_MONITOR_LANE_WIDTH_const_net_6  = 3'h0;
assign TX_DATA_2_const_net_5               = 4'h0;
assign TX_DATA_3_const_net_5               = 4'h0;
assign TX_DATA_4_const_net_5               = 4'h0;
assign TX_DATA_5_const_net_5               = 4'h0;
assign TX_DATA_6_const_net_5               = 4'h0;
assign TX_DATA_7_const_net_5               = 4'h0;
assign TX_DATA_8_const_net_5               = 4'h0;
assign TX_DATA_9_const_net_5               = 4'h0;
assign TX_DATA_10_const_net_5              = 4'h0;
assign TX_DATA_11_const_net_5              = 4'h0;
assign TX_DATA_12_const_net_6              = 4'h0;
assign TX_DATA_13_const_net_6              = 4'h0;
assign TX_DATA_14_const_net_6              = 4'h0;
assign TX_DATA_15_const_net_6              = 4'h0;
assign TX_DATA_16_const_net_6              = 4'h0;
assign TX_DATA_17_const_net_6              = 4'h0;
assign TX_DATA_18_const_net_6              = 4'h0;
assign TX_DATA_19_const_net_6              = 4'h0;
assign TX_DATA_20_const_net_6              = 4'h0;
assign TX_DATA_21_const_net_6              = 4'h0;
assign TX_DATA_22_const_net_6              = 4'h0;
assign TX_DATA_23_const_net_6              = 4'h0;
assign TX_DATA_24_const_net_6              = 4'h0;
assign TX_DATA_25_const_net_6              = 4'h0;
assign TX_DATA_26_const_net_6              = 4'h0;
assign TX_DATA_27_const_net_6              = 4'h0;
assign TX_DATA_28_const_net_6              = 4'h0;
assign TX_DATA_29_const_net_6              = 4'h0;
assign TX_DATA_30_const_net_6              = 4'h0;
assign TX_DATA_31_const_net_6              = 4'h0;
assign TX_DATA_32_const_net_6              = 4'h0;
assign TX_DATA_33_const_net_6              = 4'h0;
assign TX_DATA_34_const_net_6              = 4'h0;
assign TX_DATA_35_const_net_6              = 4'h0;
assign TX_DATA_36_const_net_6              = 4'h0;
assign TX_DATA_37_const_net_6              = 4'h0;
assign TX_DATA_38_const_net_6              = 4'h0;
assign TX_DATA_39_const_net_6              = 4'h0;
assign TX_DATA_40_const_net_6              = 4'h0;
assign TX_DATA_41_const_net_6              = 4'h0;
assign TX_DATA_42_const_net_6              = 4'h0;
assign TX_DATA_43_const_net_6              = 4'h0;
assign TX_DATA_44_const_net_6              = 4'h0;
assign TX_DATA_45_const_net_6              = 4'h0;
assign TX_DATA_46_const_net_6              = 4'h0;
assign TX_DATA_47_const_net_6              = 4'h0;
assign TX_DATA_48_const_net_6              = 4'h0;
assign TX_DATA_49_const_net_6              = 4'h0;
assign TX_DATA_50_const_net_6              = 4'h0;
assign TX_DATA_51_const_net_6              = 4'h0;
assign TX_DATA_52_const_net_6              = 4'h0;
assign TX_DATA_53_const_net_6              = 4'h0;
assign TX_DATA_54_const_net_6              = 4'h0;
assign TX_DATA_55_const_net_6              = 4'h0;
assign TX_DATA_56_const_net_6              = 4'h0;
assign TX_DATA_57_const_net_6              = 4'h0;
assign TX_DATA_58_const_net_6              = 4'h0;
assign TX_DATA_59_const_net_6              = 4'h0;
assign TX_DATA_60_const_net_6              = 4'h0;
assign TX_DATA_61_const_net_6              = 4'h0;
assign TX_DATA_62_const_net_6              = 4'h0;
assign TX_DATA_63_const_net_6              = 4'h0;
assign TX_DATA_64_const_net_6              = 4'h0;
assign TX_DATA_65_const_net_6              = 4'h0;
assign TX_DATA_66_const_net_6              = 4'h0;
assign TX_DATA_67_const_net_6              = 4'h0;
assign TX_DATA_68_const_net_6              = 4'h0;
assign TX_DATA_69_const_net_6              = 4'h0;
assign TX_DATA_70_const_net_6              = 4'h0;
assign TX_DATA_71_const_net_6              = 4'h0;
assign TX_DATA_72_const_net_6              = 4'h0;
assign TX_DATA_73_const_net_6              = 4'h0;
assign TX_DATA_74_const_net_6              = 4'h0;
assign TX_DATA_75_const_net_6              = 4'h0;
assign TX_DATA_76_const_net_6              = 4'h0;
assign TX_DATA_77_const_net_6              = 4'h0;
assign TX_DATA_78_const_net_6              = 4'h0;
assign TX_DATA_79_const_net_6              = 4'h0;
assign TX_DATA_80_const_net_6              = 4'h0;
assign TX_DATA_81_const_net_6              = 4'h0;
assign TX_DATA_82_const_net_6              = 4'h0;
assign TX_DATA_83_const_net_6              = 4'h0;
assign TX_DATA_84_const_net_6              = 4'h0;
assign TX_DATA_85_const_net_6              = 4'h0;
assign TX_DATA_86_const_net_6              = 4'h0;
assign TX_DATA_87_const_net_6              = 4'h0;
assign TX_DATA_88_const_net_6              = 4'h0;
assign TX_DATA_89_const_net_6              = 4'h0;
assign TX_DATA_90_const_net_6              = 4'h0;
assign TX_DATA_91_const_net_6              = 4'h0;
assign TX_DATA_92_const_net_6              = 4'h0;
assign TX_DATA_93_const_net_6              = 4'h0;
assign TX_DATA_94_const_net_6              = 4'h0;
assign TX_DATA_95_const_net_6              = 4'h0;
assign TX_DATA_96_const_net_6              = 4'h0;
assign TX_DATA_97_const_net_6              = 4'h0;
assign TX_DATA_98_const_net_6              = 4'h0;
assign TX_DATA_99_const_net_6              = 4'h0;
assign TX_DATA_100_const_net_6             = 4'h0;
assign TX_DATA_101_const_net_6             = 4'h0;
assign TX_DATA_102_const_net_6             = 4'h0;
assign TX_DATA_103_const_net_6             = 4'h0;
assign TX_DATA_104_const_net_6             = 4'h0;
assign TX_DATA_105_const_net_6             = 4'h0;
assign TX_DATA_106_const_net_6             = 4'h0;
assign TX_DATA_107_const_net_6             = 4'h0;
assign TX_DATA_108_const_net_6             = 4'h0;
assign TX_DATA_109_const_net_6             = 4'h0;
assign TX_DATA_110_const_net_6             = 4'h0;
assign TX_DATA_111_const_net_6             = 4'h0;
assign TX_DATA_112_const_net_6             = 4'h0;
assign TX_DATA_113_const_net_6             = 4'h0;
assign TX_DATA_114_const_net_6             = 4'h0;
assign TX_DATA_115_const_net_6             = 4'h0;
assign TX_DATA_116_const_net_6             = 4'h0;
assign TX_DATA_117_const_net_6             = 4'h0;
assign TX_DATA_118_const_net_6             = 4'h0;
assign TX_DATA_119_const_net_6             = 4'h0;
assign TX_DATA_120_const_net_6             = 4'h0;
assign TX_DATA_121_const_net_6             = 4'h0;
assign TX_DATA_122_const_net_6             = 4'h0;
assign TX_DATA_123_const_net_6             = 4'h0;
assign TX_DATA_124_const_net_6             = 4'h0;
assign TX_DATA_125_const_net_6             = 4'h0;
assign TX_DATA_126_const_net_6             = 4'h0;
assign TX_DATA_127_const_net_6             = 4'h0;
assign OE_DATA_2_const_net_6               = 4'h0;
assign OE_DATA_3_const_net_6               = 4'h0;
assign OE_DATA_4_const_net_6               = 4'h0;
assign OE_DATA_5_const_net_6               = 4'h0;
assign OE_DATA_6_const_net_6               = 4'h0;
assign OE_DATA_7_const_net_6               = 4'h0;
assign OE_DATA_8_const_net_6               = 4'h0;
assign OE_DATA_9_const_net_6               = 4'h0;
assign OE_DATA_10_const_net_6              = 4'h0;
assign OE_DATA_11_const_net_6              = 4'h0;
assign OE_DATA_12_const_net_6              = 4'h0;
assign OE_DATA_13_const_net_6              = 4'h0;
assign OE_DATA_14_const_net_6              = 4'h0;
assign OE_DATA_15_const_net_6              = 4'h0;
assign OE_DATA_16_const_net_6              = 4'h0;
assign OE_DATA_17_const_net_6              = 4'h0;
assign OE_DATA_18_const_net_6              = 4'h0;
assign OE_DATA_19_const_net_6              = 4'h0;
assign OE_DATA_20_const_net_6              = 4'h0;
assign OE_DATA_21_const_net_6              = 4'h0;
assign OE_DATA_22_const_net_6              = 4'h0;
assign OE_DATA_23_const_net_6              = 4'h0;
assign OE_DATA_24_const_net_6              = 4'h0;
assign OE_DATA_25_const_net_6              = 4'h0;
assign OE_DATA_26_const_net_6              = 4'h0;
assign OE_DATA_27_const_net_6              = 4'h0;
assign OE_DATA_28_const_net_6              = 4'h0;
assign OE_DATA_29_const_net_6              = 4'h0;
assign OE_DATA_30_const_net_6              = 4'h0;
assign OE_DATA_31_const_net_6              = 4'h0;
assign OE_DATA_32_const_net_6              = 4'h0;
assign OE_DATA_33_const_net_6              = 4'h0;
assign OE_DATA_34_const_net_6              = 4'h0;
assign OE_DATA_35_const_net_6              = 4'h0;
assign OE_DATA_36_const_net_6              = 4'h0;
assign OE_DATA_37_const_net_6              = 4'h0;
assign OE_DATA_38_const_net_6              = 4'h0;
assign OE_DATA_39_const_net_6              = 4'h0;
assign OE_DATA_40_const_net_6              = 4'h0;
assign OE_DATA_41_const_net_6              = 4'h0;
assign OE_DATA_42_const_net_6              = 4'h0;
assign OE_DATA_43_const_net_6              = 4'h0;
assign OE_DATA_44_const_net_6              = 4'h0;
assign OE_DATA_45_const_net_6              = 4'h0;
assign OE_DATA_46_const_net_6              = 4'h0;
assign OE_DATA_47_const_net_6              = 4'h0;
assign OE_DATA_48_const_net_6              = 4'h0;
assign OE_DATA_49_const_net_6              = 4'h0;
assign OE_DATA_50_const_net_6              = 4'h0;
assign OE_DATA_51_const_net_6              = 4'h0;
assign OE_DATA_52_const_net_6              = 4'h0;
assign OE_DATA_53_const_net_6              = 4'h0;
assign OE_DATA_54_const_net_6              = 4'h0;
assign OE_DATA_55_const_net_6              = 4'h0;
assign OE_DATA_56_const_net_6              = 4'h0;
assign OE_DATA_57_const_net_6              = 4'h0;
assign OE_DATA_58_const_net_6              = 4'h0;
assign OE_DATA_59_const_net_6              = 4'h0;
assign OE_DATA_60_const_net_6              = 4'h0;
assign OE_DATA_61_const_net_6              = 4'h0;
assign OE_DATA_62_const_net_6              = 4'h0;
assign OE_DATA_63_const_net_6              = 4'h0;
assign OE_DATA_64_const_net_6              = 4'h0;
assign OE_DATA_65_const_net_6              = 4'h0;
assign OE_DATA_66_const_net_6              = 4'h0;
assign OE_DATA_67_const_net_6              = 4'h0;
assign OE_DATA_68_const_net_6              = 4'h0;
assign OE_DATA_69_const_net_6              = 4'h0;
assign OE_DATA_70_const_net_6              = 4'h0;
assign OE_DATA_71_const_net_6              = 4'h0;
assign OE_DATA_72_const_net_6              = 4'h0;
assign OE_DATA_73_const_net_6              = 4'h0;
assign OE_DATA_74_const_net_6              = 4'h0;
assign OE_DATA_75_const_net_6              = 4'h0;
assign OE_DATA_76_const_net_6              = 4'h0;
assign OE_DATA_77_const_net_6              = 4'h0;
assign OE_DATA_78_const_net_6              = 4'h0;
assign OE_DATA_79_const_net_6              = 4'h0;
assign OE_DATA_80_const_net_6              = 4'h0;
assign OE_DATA_81_const_net_6              = 4'h0;
assign OE_DATA_82_const_net_6              = 4'h0;
assign OE_DATA_83_const_net_6              = 4'h0;
assign OE_DATA_84_const_net_6              = 4'h0;
assign OE_DATA_85_const_net_6              = 4'h0;
assign OE_DATA_86_const_net_6              = 4'h0;
assign OE_DATA_87_const_net_6              = 4'h0;
assign OE_DATA_88_const_net_6              = 4'h0;
assign OE_DATA_89_const_net_6              = 4'h0;
assign OE_DATA_90_const_net_6              = 4'h0;
assign OE_DATA_91_const_net_6              = 4'h0;
assign OE_DATA_92_const_net_6              = 4'h0;
assign OE_DATA_93_const_net_6              = 4'h0;
assign OE_DATA_94_const_net_6              = 4'h0;
assign OE_DATA_95_const_net_6              = 4'h0;
assign OE_DATA_96_const_net_6              = 4'h0;
assign OE_DATA_97_const_net_6              = 4'h0;
assign OE_DATA_98_const_net_6              = 4'h0;
assign OE_DATA_99_const_net_6              = 4'h0;
assign OE_DATA_100_const_net_6             = 4'h0;
assign OE_DATA_101_const_net_6             = 4'h0;
assign OE_DATA_102_const_net_6             = 4'h0;
assign OE_DATA_103_const_net_6             = 4'h0;
assign OE_DATA_104_const_net_6             = 4'h0;
assign OE_DATA_105_const_net_6             = 4'h0;
assign OE_DATA_106_const_net_6             = 4'h0;
assign OE_DATA_107_const_net_6             = 4'h0;
assign OE_DATA_108_const_net_6             = 4'h0;
assign OE_DATA_109_const_net_6             = 4'h0;
assign OE_DATA_110_const_net_6             = 4'h0;
assign OE_DATA_111_const_net_6             = 4'h0;
assign OE_DATA_112_const_net_6             = 4'h0;
assign OE_DATA_113_const_net_6             = 4'h0;
assign OE_DATA_114_const_net_6             = 4'h0;
assign OE_DATA_115_const_net_6             = 4'h0;
assign OE_DATA_116_const_net_6             = 4'h0;
assign OE_DATA_117_const_net_6             = 4'h0;
assign OE_DATA_118_const_net_6             = 4'h0;
assign OE_DATA_119_const_net_6             = 4'h0;
assign OE_DATA_120_const_net_6             = 4'h0;
assign OE_DATA_121_const_net_6             = 4'h0;
assign OE_DATA_122_const_net_6             = 4'h0;
assign OE_DATA_123_const_net_6             = 4'h0;
assign OE_DATA_124_const_net_6             = 4'h0;
assign OE_DATA_125_const_net_6             = 4'h0;
assign OE_DATA_126_const_net_6             = 4'h0;
assign OE_DATA_127_const_net_6             = 4'h0;
assign PAD_const_net_2                     = 2'h0;
assign PAD_I_const_net_2                   = 2'h0;
assign PAD_N_const_net_2                   = 2'h0;
assign PAD_I_N_const_net_2                 = 2'h0;
assign RX_DQS_90_const_net_7               = 2'h0;
assign FIFO_WR_PTR_const_net_7             = 3'h0;
assign FIFO_RD_PTR_const_net_7             = 3'h0;
assign EYE_MONITOR_LANE_WIDTH_const_net_7  = 3'h0;
assign TX_DATA_1_const_net_4               = 4'h0;
assign TX_DATA_2_const_net_6               = 4'h0;
assign TX_DATA_3_const_net_6               = 4'h0;
assign TX_DATA_4_const_net_6               = 4'h0;
assign TX_DATA_5_const_net_6               = 4'h0;
assign TX_DATA_6_const_net_6               = 4'h0;
assign TX_DATA_7_const_net_6               = 4'h0;
assign TX_DATA_8_const_net_6               = 4'h0;
assign TX_DATA_9_const_net_6               = 4'h0;
assign TX_DATA_10_const_net_6              = 4'h0;
assign TX_DATA_11_const_net_6              = 4'h0;
assign TX_DATA_12_const_net_7              = 4'h0;
assign TX_DATA_13_const_net_7              = 4'h0;
assign TX_DATA_14_const_net_7              = 4'h0;
assign TX_DATA_15_const_net_7              = 4'h0;
assign TX_DATA_16_const_net_7              = 4'h0;
assign TX_DATA_17_const_net_7              = 4'h0;
assign TX_DATA_18_const_net_7              = 4'h0;
assign TX_DATA_19_const_net_7              = 4'h0;
assign TX_DATA_20_const_net_7              = 4'h0;
assign TX_DATA_21_const_net_7              = 4'h0;
assign TX_DATA_22_const_net_7              = 4'h0;
assign TX_DATA_23_const_net_7              = 4'h0;
assign TX_DATA_24_const_net_7              = 4'h0;
assign TX_DATA_25_const_net_7              = 4'h0;
assign TX_DATA_26_const_net_7              = 4'h0;
assign TX_DATA_27_const_net_7              = 4'h0;
assign TX_DATA_28_const_net_7              = 4'h0;
assign TX_DATA_29_const_net_7              = 4'h0;
assign TX_DATA_30_const_net_7              = 4'h0;
assign TX_DATA_31_const_net_7              = 4'h0;
assign TX_DATA_32_const_net_7              = 4'h0;
assign TX_DATA_33_const_net_7              = 4'h0;
assign TX_DATA_34_const_net_7              = 4'h0;
assign TX_DATA_35_const_net_7              = 4'h0;
assign TX_DATA_36_const_net_7              = 4'h0;
assign TX_DATA_37_const_net_7              = 4'h0;
assign TX_DATA_38_const_net_7              = 4'h0;
assign TX_DATA_39_const_net_7              = 4'h0;
assign TX_DATA_40_const_net_7              = 4'h0;
assign TX_DATA_41_const_net_7              = 4'h0;
assign TX_DATA_42_const_net_7              = 4'h0;
assign TX_DATA_43_const_net_7              = 4'h0;
assign TX_DATA_44_const_net_7              = 4'h0;
assign TX_DATA_45_const_net_7              = 4'h0;
assign TX_DATA_46_const_net_7              = 4'h0;
assign TX_DATA_47_const_net_7              = 4'h0;
assign TX_DATA_48_const_net_7              = 4'h0;
assign TX_DATA_49_const_net_7              = 4'h0;
assign TX_DATA_50_const_net_7              = 4'h0;
assign TX_DATA_51_const_net_7              = 4'h0;
assign TX_DATA_52_const_net_7              = 4'h0;
assign TX_DATA_53_const_net_7              = 4'h0;
assign TX_DATA_54_const_net_7              = 4'h0;
assign TX_DATA_55_const_net_7              = 4'h0;
assign TX_DATA_56_const_net_7              = 4'h0;
assign TX_DATA_57_const_net_7              = 4'h0;
assign TX_DATA_58_const_net_7              = 4'h0;
assign TX_DATA_59_const_net_7              = 4'h0;
assign TX_DATA_60_const_net_7              = 4'h0;
assign TX_DATA_61_const_net_7              = 4'h0;
assign TX_DATA_62_const_net_7              = 4'h0;
assign TX_DATA_63_const_net_7              = 4'h0;
assign TX_DATA_64_const_net_7              = 4'h0;
assign TX_DATA_65_const_net_7              = 4'h0;
assign TX_DATA_66_const_net_7              = 4'h0;
assign TX_DATA_67_const_net_7              = 4'h0;
assign TX_DATA_68_const_net_7              = 4'h0;
assign TX_DATA_69_const_net_7              = 4'h0;
assign TX_DATA_70_const_net_7              = 4'h0;
assign TX_DATA_71_const_net_7              = 4'h0;
assign TX_DATA_72_const_net_7              = 4'h0;
assign TX_DATA_73_const_net_7              = 4'h0;
assign TX_DATA_74_const_net_7              = 4'h0;
assign TX_DATA_75_const_net_7              = 4'h0;
assign TX_DATA_76_const_net_7              = 4'h0;
assign TX_DATA_77_const_net_7              = 4'h0;
assign TX_DATA_78_const_net_7              = 4'h0;
assign TX_DATA_79_const_net_7              = 4'h0;
assign TX_DATA_80_const_net_7              = 4'h0;
assign TX_DATA_81_const_net_7              = 4'h0;
assign TX_DATA_82_const_net_7              = 4'h0;
assign TX_DATA_83_const_net_7              = 4'h0;
assign TX_DATA_84_const_net_7              = 4'h0;
assign TX_DATA_85_const_net_7              = 4'h0;
assign TX_DATA_86_const_net_7              = 4'h0;
assign TX_DATA_87_const_net_7              = 4'h0;
assign TX_DATA_88_const_net_7              = 4'h0;
assign TX_DATA_89_const_net_7              = 4'h0;
assign TX_DATA_90_const_net_7              = 4'h0;
assign TX_DATA_91_const_net_7              = 4'h0;
assign TX_DATA_92_const_net_7              = 4'h0;
assign TX_DATA_93_const_net_7              = 4'h0;
assign TX_DATA_94_const_net_7              = 4'h0;
assign TX_DATA_95_const_net_7              = 4'h0;
assign TX_DATA_96_const_net_7              = 4'h0;
assign TX_DATA_97_const_net_7              = 4'h0;
assign TX_DATA_98_const_net_7              = 4'h0;
assign TX_DATA_99_const_net_7              = 4'h0;
assign TX_DATA_100_const_net_7             = 4'h0;
assign TX_DATA_101_const_net_7             = 4'h0;
assign TX_DATA_102_const_net_7             = 4'h0;
assign TX_DATA_103_const_net_7             = 4'h0;
assign TX_DATA_104_const_net_7             = 4'h0;
assign TX_DATA_105_const_net_7             = 4'h0;
assign TX_DATA_106_const_net_7             = 4'h0;
assign TX_DATA_107_const_net_7             = 4'h0;
assign TX_DATA_108_const_net_7             = 4'h0;
assign TX_DATA_109_const_net_7             = 4'h0;
assign TX_DATA_110_const_net_7             = 4'h0;
assign TX_DATA_111_const_net_7             = 4'h0;
assign TX_DATA_112_const_net_7             = 4'h0;
assign TX_DATA_113_const_net_7             = 4'h0;
assign TX_DATA_114_const_net_7             = 4'h0;
assign TX_DATA_115_const_net_7             = 4'h0;
assign TX_DATA_116_const_net_7             = 4'h0;
assign TX_DATA_117_const_net_7             = 4'h0;
assign TX_DATA_118_const_net_7             = 4'h0;
assign TX_DATA_119_const_net_7             = 4'h0;
assign TX_DATA_120_const_net_7             = 4'h0;
assign TX_DATA_121_const_net_7             = 4'h0;
assign TX_DATA_122_const_net_7             = 4'h0;
assign TX_DATA_123_const_net_7             = 4'h0;
assign TX_DATA_124_const_net_7             = 4'h0;
assign TX_DATA_125_const_net_7             = 4'h0;
assign TX_DATA_126_const_net_7             = 4'h0;
assign TX_DATA_127_const_net_7             = 4'h0;
assign OE_DATA_1_const_net_7               = 4'h0;
assign OE_DATA_2_const_net_7               = 4'h0;
assign OE_DATA_3_const_net_7               = 4'h0;
assign OE_DATA_4_const_net_7               = 4'h0;
assign OE_DATA_5_const_net_7               = 4'h0;
assign OE_DATA_6_const_net_7               = 4'h0;
assign OE_DATA_7_const_net_7               = 4'h0;
assign OE_DATA_8_const_net_7               = 4'h0;
assign OE_DATA_9_const_net_7               = 4'h0;
assign OE_DATA_10_const_net_7              = 4'h0;
assign OE_DATA_11_const_net_7              = 4'h0;
assign OE_DATA_12_const_net_7              = 4'h0;
assign OE_DATA_13_const_net_7              = 4'h0;
assign OE_DATA_14_const_net_7              = 4'h0;
assign OE_DATA_15_const_net_7              = 4'h0;
assign OE_DATA_16_const_net_7              = 4'h0;
assign OE_DATA_17_const_net_7              = 4'h0;
assign OE_DATA_18_const_net_7              = 4'h0;
assign OE_DATA_19_const_net_7              = 4'h0;
assign OE_DATA_20_const_net_7              = 4'h0;
assign OE_DATA_21_const_net_7              = 4'h0;
assign OE_DATA_22_const_net_7              = 4'h0;
assign OE_DATA_23_const_net_7              = 4'h0;
assign OE_DATA_24_const_net_7              = 4'h0;
assign OE_DATA_25_const_net_7              = 4'h0;
assign OE_DATA_26_const_net_7              = 4'h0;
assign OE_DATA_27_const_net_7              = 4'h0;
assign OE_DATA_28_const_net_7              = 4'h0;
assign OE_DATA_29_const_net_7              = 4'h0;
assign OE_DATA_30_const_net_7              = 4'h0;
assign OE_DATA_31_const_net_7              = 4'h0;
assign OE_DATA_32_const_net_7              = 4'h0;
assign OE_DATA_33_const_net_7              = 4'h0;
assign OE_DATA_34_const_net_7              = 4'h0;
assign OE_DATA_35_const_net_7              = 4'h0;
assign OE_DATA_36_const_net_7              = 4'h0;
assign OE_DATA_37_const_net_7              = 4'h0;
assign OE_DATA_38_const_net_7              = 4'h0;
assign OE_DATA_39_const_net_7              = 4'h0;
assign OE_DATA_40_const_net_7              = 4'h0;
assign OE_DATA_41_const_net_7              = 4'h0;
assign OE_DATA_42_const_net_7              = 4'h0;
assign OE_DATA_43_const_net_7              = 4'h0;
assign OE_DATA_44_const_net_7              = 4'h0;
assign OE_DATA_45_const_net_7              = 4'h0;
assign OE_DATA_46_const_net_7              = 4'h0;
assign OE_DATA_47_const_net_7              = 4'h0;
assign OE_DATA_48_const_net_7              = 4'h0;
assign OE_DATA_49_const_net_7              = 4'h0;
assign OE_DATA_50_const_net_7              = 4'h0;
assign OE_DATA_51_const_net_7              = 4'h0;
assign OE_DATA_52_const_net_7              = 4'h0;
assign OE_DATA_53_const_net_7              = 4'h0;
assign OE_DATA_54_const_net_7              = 4'h0;
assign OE_DATA_55_const_net_7              = 4'h0;
assign OE_DATA_56_const_net_7              = 4'h0;
assign OE_DATA_57_const_net_7              = 4'h0;
assign OE_DATA_58_const_net_7              = 4'h0;
assign OE_DATA_59_const_net_7              = 4'h0;
assign OE_DATA_60_const_net_7              = 4'h0;
assign OE_DATA_61_const_net_7              = 4'h0;
assign OE_DATA_62_const_net_7              = 4'h0;
assign OE_DATA_63_const_net_7              = 4'h0;
assign OE_DATA_64_const_net_7              = 4'h0;
assign OE_DATA_65_const_net_7              = 4'h0;
assign OE_DATA_66_const_net_7              = 4'h0;
assign OE_DATA_67_const_net_7              = 4'h0;
assign OE_DATA_68_const_net_7              = 4'h0;
assign OE_DATA_69_const_net_7              = 4'h0;
assign OE_DATA_70_const_net_7              = 4'h0;
assign OE_DATA_71_const_net_7              = 4'h0;
assign OE_DATA_72_const_net_7              = 4'h0;
assign OE_DATA_73_const_net_7              = 4'h0;
assign OE_DATA_74_const_net_7              = 4'h0;
assign OE_DATA_75_const_net_7              = 4'h0;
assign OE_DATA_76_const_net_7              = 4'h0;
assign OE_DATA_77_const_net_7              = 4'h0;
assign OE_DATA_78_const_net_7              = 4'h0;
assign OE_DATA_79_const_net_7              = 4'h0;
assign OE_DATA_80_const_net_7              = 4'h0;
assign OE_DATA_81_const_net_7              = 4'h0;
assign OE_DATA_82_const_net_7              = 4'h0;
assign OE_DATA_83_const_net_7              = 4'h0;
assign OE_DATA_84_const_net_7              = 4'h0;
assign OE_DATA_85_const_net_7              = 4'h0;
assign OE_DATA_86_const_net_7              = 4'h0;
assign OE_DATA_87_const_net_7              = 4'h0;
assign OE_DATA_88_const_net_7              = 4'h0;
assign OE_DATA_89_const_net_7              = 4'h0;
assign OE_DATA_90_const_net_7              = 4'h0;
assign OE_DATA_91_const_net_7              = 4'h0;
assign OE_DATA_92_const_net_7              = 4'h0;
assign OE_DATA_93_const_net_7              = 4'h0;
assign OE_DATA_94_const_net_7              = 4'h0;
assign OE_DATA_95_const_net_7              = 4'h0;
assign OE_DATA_96_const_net_7              = 4'h0;
assign OE_DATA_97_const_net_7              = 4'h0;
assign OE_DATA_98_const_net_7              = 4'h0;
assign OE_DATA_99_const_net_7              = 4'h0;
assign OE_DATA_100_const_net_7             = 4'h0;
assign OE_DATA_101_const_net_7             = 4'h0;
assign OE_DATA_102_const_net_7             = 4'h0;
assign OE_DATA_103_const_net_7             = 4'h0;
assign OE_DATA_104_const_net_7             = 4'h0;
assign OE_DATA_105_const_net_7             = 4'h0;
assign OE_DATA_106_const_net_7             = 4'h0;
assign OE_DATA_107_const_net_7             = 4'h0;
assign OE_DATA_108_const_net_7             = 4'h0;
assign OE_DATA_109_const_net_7             = 4'h0;
assign OE_DATA_110_const_net_7             = 4'h0;
assign OE_DATA_111_const_net_7             = 4'h0;
assign OE_DATA_112_const_net_7             = 4'h0;
assign OE_DATA_113_const_net_7             = 4'h0;
assign OE_DATA_114_const_net_7             = 4'h0;
assign OE_DATA_115_const_net_7             = 4'h0;
assign OE_DATA_116_const_net_7             = 4'h0;
assign OE_DATA_117_const_net_7             = 4'h0;
assign OE_DATA_118_const_net_7             = 4'h0;
assign OE_DATA_119_const_net_7             = 4'h0;
assign OE_DATA_120_const_net_7             = 4'h0;
assign OE_DATA_121_const_net_7             = 4'h0;
assign OE_DATA_122_const_net_7             = 4'h0;
assign OE_DATA_123_const_net_7             = 4'h0;
assign OE_DATA_124_const_net_7             = 4'h0;
assign OE_DATA_125_const_net_7             = 4'h0;
assign OE_DATA_126_const_net_7             = 4'h0;
assign OE_DATA_127_const_net_7             = 4'h0;
assign RX_DQS_90_const_net_8               = 2'h0;
assign FIFO_WR_PTR_const_net_8             = 3'h0;
assign FIFO_RD_PTR_const_net_8             = 3'h0;
assign EYE_MONITOR_LANE_WIDTH_const_net_8  = 3'h0;
assign TX_DATA_1_const_net_5               = 4'h0;
assign TX_DATA_2_const_net_7               = 4'h0;
assign TX_DATA_3_const_net_7               = 4'h0;
assign TX_DATA_4_const_net_7               = 4'h0;
assign TX_DATA_5_const_net_7               = 4'h0;
assign TX_DATA_6_const_net_7               = 4'h0;
assign TX_DATA_7_const_net_7               = 4'h0;
assign TX_DATA_8_const_net_7               = 4'h0;
assign TX_DATA_9_const_net_7               = 4'h0;
assign TX_DATA_10_const_net_7              = 4'h0;
assign TX_DATA_11_const_net_7              = 4'h0;
assign TX_DATA_12_const_net_8              = 4'h0;
assign TX_DATA_13_const_net_8              = 4'h0;
assign TX_DATA_14_const_net_8              = 4'h0;
assign TX_DATA_15_const_net_8              = 4'h0;
assign TX_DATA_16_const_net_8              = 4'h0;
assign TX_DATA_17_const_net_8              = 4'h0;
assign TX_DATA_18_const_net_8              = 4'h0;
assign TX_DATA_19_const_net_8              = 4'h0;
assign TX_DATA_20_const_net_8              = 4'h0;
assign TX_DATA_21_const_net_8              = 4'h0;
assign TX_DATA_22_const_net_8              = 4'h0;
assign TX_DATA_23_const_net_8              = 4'h0;
assign TX_DATA_24_const_net_8              = 4'h0;
assign TX_DATA_25_const_net_8              = 4'h0;
assign TX_DATA_26_const_net_8              = 4'h0;
assign TX_DATA_27_const_net_8              = 4'h0;
assign TX_DATA_28_const_net_8              = 4'h0;
assign TX_DATA_29_const_net_8              = 4'h0;
assign TX_DATA_30_const_net_8              = 4'h0;
assign TX_DATA_31_const_net_8              = 4'h0;
assign TX_DATA_32_const_net_8              = 4'h0;
assign TX_DATA_33_const_net_8              = 4'h0;
assign TX_DATA_34_const_net_8              = 4'h0;
assign TX_DATA_35_const_net_8              = 4'h0;
assign TX_DATA_36_const_net_8              = 4'h0;
assign TX_DATA_37_const_net_8              = 4'h0;
assign TX_DATA_38_const_net_8              = 4'h0;
assign TX_DATA_39_const_net_8              = 4'h0;
assign TX_DATA_40_const_net_8              = 4'h0;
assign TX_DATA_41_const_net_8              = 4'h0;
assign TX_DATA_42_const_net_8              = 4'h0;
assign TX_DATA_43_const_net_8              = 4'h0;
assign TX_DATA_44_const_net_8              = 4'h0;
assign TX_DATA_45_const_net_8              = 4'h0;
assign TX_DATA_46_const_net_8              = 4'h0;
assign TX_DATA_47_const_net_8              = 4'h0;
assign TX_DATA_48_const_net_8              = 4'h0;
assign TX_DATA_49_const_net_8              = 4'h0;
assign TX_DATA_50_const_net_8              = 4'h0;
assign TX_DATA_51_const_net_8              = 4'h0;
assign TX_DATA_52_const_net_8              = 4'h0;
assign TX_DATA_53_const_net_8              = 4'h0;
assign TX_DATA_54_const_net_8              = 4'h0;
assign TX_DATA_55_const_net_8              = 4'h0;
assign TX_DATA_56_const_net_8              = 4'h0;
assign TX_DATA_57_const_net_8              = 4'h0;
assign TX_DATA_58_const_net_8              = 4'h0;
assign TX_DATA_59_const_net_8              = 4'h0;
assign TX_DATA_60_const_net_8              = 4'h0;
assign TX_DATA_61_const_net_8              = 4'h0;
assign TX_DATA_62_const_net_8              = 4'h0;
assign TX_DATA_63_const_net_8              = 4'h0;
assign TX_DATA_64_const_net_8              = 4'h0;
assign TX_DATA_65_const_net_8              = 4'h0;
assign TX_DATA_66_const_net_8              = 4'h0;
assign TX_DATA_67_const_net_8              = 4'h0;
assign TX_DATA_68_const_net_8              = 4'h0;
assign TX_DATA_69_const_net_8              = 4'h0;
assign TX_DATA_70_const_net_8              = 4'h0;
assign TX_DATA_71_const_net_8              = 4'h0;
assign TX_DATA_72_const_net_8              = 4'h0;
assign TX_DATA_73_const_net_8              = 4'h0;
assign TX_DATA_74_const_net_8              = 4'h0;
assign TX_DATA_75_const_net_8              = 4'h0;
assign TX_DATA_76_const_net_8              = 4'h0;
assign TX_DATA_77_const_net_8              = 4'h0;
assign TX_DATA_78_const_net_8              = 4'h0;
assign TX_DATA_79_const_net_8              = 4'h0;
assign TX_DATA_80_const_net_8              = 4'h0;
assign TX_DATA_81_const_net_8              = 4'h0;
assign TX_DATA_82_const_net_8              = 4'h0;
assign TX_DATA_83_const_net_8              = 4'h0;
assign TX_DATA_84_const_net_8              = 4'h0;
assign TX_DATA_85_const_net_8              = 4'h0;
assign TX_DATA_86_const_net_8              = 4'h0;
assign TX_DATA_87_const_net_8              = 4'h0;
assign TX_DATA_88_const_net_8              = 4'h0;
assign TX_DATA_89_const_net_8              = 4'h0;
assign TX_DATA_90_const_net_8              = 4'h0;
assign TX_DATA_91_const_net_8              = 4'h0;
assign TX_DATA_92_const_net_8              = 4'h0;
assign TX_DATA_93_const_net_8              = 4'h0;
assign TX_DATA_94_const_net_8              = 4'h0;
assign TX_DATA_95_const_net_8              = 4'h0;
assign TX_DATA_96_const_net_8              = 4'h0;
assign TX_DATA_97_const_net_8              = 4'h0;
assign TX_DATA_98_const_net_8              = 4'h0;
assign TX_DATA_99_const_net_8              = 4'h0;
assign TX_DATA_100_const_net_8             = 4'h0;
assign TX_DATA_101_const_net_8             = 4'h0;
assign TX_DATA_102_const_net_8             = 4'h0;
assign TX_DATA_103_const_net_8             = 4'h0;
assign TX_DATA_104_const_net_8             = 4'h0;
assign TX_DATA_105_const_net_8             = 4'h0;
assign TX_DATA_106_const_net_8             = 4'h0;
assign TX_DATA_107_const_net_8             = 4'h0;
assign TX_DATA_108_const_net_8             = 4'h0;
assign TX_DATA_109_const_net_8             = 4'h0;
assign TX_DATA_110_const_net_8             = 4'h0;
assign TX_DATA_111_const_net_8             = 4'h0;
assign TX_DATA_112_const_net_8             = 4'h0;
assign TX_DATA_113_const_net_8             = 4'h0;
assign TX_DATA_114_const_net_8             = 4'h0;
assign TX_DATA_115_const_net_8             = 4'h0;
assign TX_DATA_116_const_net_8             = 4'h0;
assign TX_DATA_117_const_net_8             = 4'h0;
assign TX_DATA_118_const_net_8             = 4'h0;
assign TX_DATA_119_const_net_8             = 4'h0;
assign TX_DATA_120_const_net_8             = 4'h0;
assign TX_DATA_121_const_net_8             = 4'h0;
assign TX_DATA_122_const_net_8             = 4'h0;
assign TX_DATA_123_const_net_8             = 4'h0;
assign TX_DATA_124_const_net_8             = 4'h0;
assign TX_DATA_125_const_net_8             = 4'h0;
assign TX_DATA_126_const_net_8             = 4'h0;
assign TX_DATA_127_const_net_8             = 4'h0;
assign OE_DATA_1_const_net_8               = 4'h0;
assign OE_DATA_2_const_net_8               = 4'h0;
assign OE_DATA_3_const_net_8               = 4'h0;
assign OE_DATA_4_const_net_8               = 4'h0;
assign OE_DATA_5_const_net_8               = 4'h0;
assign OE_DATA_6_const_net_8               = 4'h0;
assign OE_DATA_7_const_net_8               = 4'h0;
assign OE_DATA_8_const_net_8               = 4'h0;
assign OE_DATA_9_const_net_8               = 4'h0;
assign OE_DATA_10_const_net_8              = 4'h0;
assign OE_DATA_11_const_net_8              = 4'h0;
assign OE_DATA_12_const_net_8              = 4'h0;
assign OE_DATA_13_const_net_8              = 4'h0;
assign OE_DATA_14_const_net_8              = 4'h0;
assign OE_DATA_15_const_net_8              = 4'h0;
assign OE_DATA_16_const_net_8              = 4'h0;
assign OE_DATA_17_const_net_8              = 4'h0;
assign OE_DATA_18_const_net_8              = 4'h0;
assign OE_DATA_19_const_net_8              = 4'h0;
assign OE_DATA_20_const_net_8              = 4'h0;
assign OE_DATA_21_const_net_8              = 4'h0;
assign OE_DATA_22_const_net_8              = 4'h0;
assign OE_DATA_23_const_net_8              = 4'h0;
assign OE_DATA_24_const_net_8              = 4'h0;
assign OE_DATA_25_const_net_8              = 4'h0;
assign OE_DATA_26_const_net_8              = 4'h0;
assign OE_DATA_27_const_net_8              = 4'h0;
assign OE_DATA_28_const_net_8              = 4'h0;
assign OE_DATA_29_const_net_8              = 4'h0;
assign OE_DATA_30_const_net_8              = 4'h0;
assign OE_DATA_31_const_net_8              = 4'h0;
assign OE_DATA_32_const_net_8              = 4'h0;
assign OE_DATA_33_const_net_8              = 4'h0;
assign OE_DATA_34_const_net_8              = 4'h0;
assign OE_DATA_35_const_net_8              = 4'h0;
assign OE_DATA_36_const_net_8              = 4'h0;
assign OE_DATA_37_const_net_8              = 4'h0;
assign OE_DATA_38_const_net_8              = 4'h0;
assign OE_DATA_39_const_net_8              = 4'h0;
assign OE_DATA_40_const_net_8              = 4'h0;
assign OE_DATA_41_const_net_8              = 4'h0;
assign OE_DATA_42_const_net_8              = 4'h0;
assign OE_DATA_43_const_net_8              = 4'h0;
assign OE_DATA_44_const_net_8              = 4'h0;
assign OE_DATA_45_const_net_8              = 4'h0;
assign OE_DATA_46_const_net_8              = 4'h0;
assign OE_DATA_47_const_net_8              = 4'h0;
assign OE_DATA_48_const_net_8              = 4'h0;
assign OE_DATA_49_const_net_8              = 4'h0;
assign OE_DATA_50_const_net_8              = 4'h0;
assign OE_DATA_51_const_net_8              = 4'h0;
assign OE_DATA_52_const_net_8              = 4'h0;
assign OE_DATA_53_const_net_8              = 4'h0;
assign OE_DATA_54_const_net_8              = 4'h0;
assign OE_DATA_55_const_net_8              = 4'h0;
assign OE_DATA_56_const_net_8              = 4'h0;
assign OE_DATA_57_const_net_8              = 4'h0;
assign OE_DATA_58_const_net_8              = 4'h0;
assign OE_DATA_59_const_net_8              = 4'h0;
assign OE_DATA_60_const_net_8              = 4'h0;
assign OE_DATA_61_const_net_8              = 4'h0;
assign OE_DATA_62_const_net_8              = 4'h0;
assign OE_DATA_63_const_net_8              = 4'h0;
assign OE_DATA_64_const_net_8              = 4'h0;
assign OE_DATA_65_const_net_8              = 4'h0;
assign OE_DATA_66_const_net_8              = 4'h0;
assign OE_DATA_67_const_net_8              = 4'h0;
assign OE_DATA_68_const_net_8              = 4'h0;
assign OE_DATA_69_const_net_8              = 4'h0;
assign OE_DATA_70_const_net_8              = 4'h0;
assign OE_DATA_71_const_net_8              = 4'h0;
assign OE_DATA_72_const_net_8              = 4'h0;
assign OE_DATA_73_const_net_8              = 4'h0;
assign OE_DATA_74_const_net_8              = 4'h0;
assign OE_DATA_75_const_net_8              = 4'h0;
assign OE_DATA_76_const_net_8              = 4'h0;
assign OE_DATA_77_const_net_8              = 4'h0;
assign OE_DATA_78_const_net_8              = 4'h0;
assign OE_DATA_79_const_net_8              = 4'h0;
assign OE_DATA_80_const_net_8              = 4'h0;
assign OE_DATA_81_const_net_8              = 4'h0;
assign OE_DATA_82_const_net_8              = 4'h0;
assign OE_DATA_83_const_net_8              = 4'h0;
assign OE_DATA_84_const_net_8              = 4'h0;
assign OE_DATA_85_const_net_8              = 4'h0;
assign OE_DATA_86_const_net_8              = 4'h0;
assign OE_DATA_87_const_net_8              = 4'h0;
assign OE_DATA_88_const_net_8              = 4'h0;
assign OE_DATA_89_const_net_8              = 4'h0;
assign OE_DATA_90_const_net_8              = 4'h0;
assign OE_DATA_91_const_net_8              = 4'h0;
assign OE_DATA_92_const_net_8              = 4'h0;
assign OE_DATA_93_const_net_8              = 4'h0;
assign OE_DATA_94_const_net_8              = 4'h0;
assign OE_DATA_95_const_net_8              = 4'h0;
assign OE_DATA_96_const_net_8              = 4'h0;
assign OE_DATA_97_const_net_8              = 4'h0;
assign OE_DATA_98_const_net_8              = 4'h0;
assign OE_DATA_99_const_net_8              = 4'h0;
assign OE_DATA_100_const_net_8             = 4'h0;
assign OE_DATA_101_const_net_8             = 4'h0;
assign OE_DATA_102_const_net_8             = 4'h0;
assign OE_DATA_103_const_net_8             = 4'h0;
assign OE_DATA_104_const_net_8             = 4'h0;
assign OE_DATA_105_const_net_8             = 4'h0;
assign OE_DATA_106_const_net_8             = 4'h0;
assign OE_DATA_107_const_net_8             = 4'h0;
assign OE_DATA_108_const_net_8             = 4'h0;
assign OE_DATA_109_const_net_8             = 4'h0;
assign OE_DATA_110_const_net_8             = 4'h0;
assign OE_DATA_111_const_net_8             = 4'h0;
assign OE_DATA_112_const_net_8             = 4'h0;
assign OE_DATA_113_const_net_8             = 4'h0;
assign OE_DATA_114_const_net_8             = 4'h0;
assign OE_DATA_115_const_net_8             = 4'h0;
assign OE_DATA_116_const_net_8             = 4'h0;
assign OE_DATA_117_const_net_8             = 4'h0;
assign OE_DATA_118_const_net_8             = 4'h0;
assign OE_DATA_119_const_net_8             = 4'h0;
assign OE_DATA_120_const_net_8             = 4'h0;
assign OE_DATA_121_const_net_8             = 4'h0;
assign OE_DATA_122_const_net_8             = 4'h0;
assign OE_DATA_123_const_net_8             = 4'h0;
assign OE_DATA_124_const_net_8             = 4'h0;
assign OE_DATA_125_const_net_8             = 4'h0;
assign OE_DATA_126_const_net_8             = 4'h0;
assign OE_DATA_127_const_net_8             = 4'h0;
assign RX_DQS_90_const_net_9               = 2'h0;
assign FIFO_WR_PTR_const_net_9             = 3'h0;
assign FIFO_RD_PTR_const_net_9             = 3'h0;
assign EYE_MONITOR_LANE_WIDTH_const_net_9  = 3'h0;
assign TX_DATA_1_const_net_6               = 4'h0;
assign TX_DATA_2_const_net_8               = 4'h0;
assign TX_DATA_3_const_net_8               = 4'h0;
assign TX_DATA_4_const_net_8               = 4'h0;
assign TX_DATA_5_const_net_8               = 4'h0;
assign TX_DATA_6_const_net_8               = 4'h0;
assign TX_DATA_7_const_net_8               = 4'h0;
assign TX_DATA_8_const_net_8               = 4'h0;
assign TX_DATA_9_const_net_8               = 4'h0;
assign TX_DATA_10_const_net_8              = 4'h0;
assign TX_DATA_11_const_net_8              = 4'h0;
assign TX_DATA_12_const_net_9              = 4'h0;
assign TX_DATA_13_const_net_9              = 4'h0;
assign TX_DATA_14_const_net_9              = 4'h0;
assign TX_DATA_15_const_net_9              = 4'h0;
assign TX_DATA_16_const_net_9              = 4'h0;
assign TX_DATA_17_const_net_9              = 4'h0;
assign TX_DATA_18_const_net_9              = 4'h0;
assign TX_DATA_19_const_net_9              = 4'h0;
assign TX_DATA_20_const_net_9              = 4'h0;
assign TX_DATA_21_const_net_9              = 4'h0;
assign TX_DATA_22_const_net_9              = 4'h0;
assign TX_DATA_23_const_net_9              = 4'h0;
assign TX_DATA_24_const_net_9              = 4'h0;
assign TX_DATA_25_const_net_9              = 4'h0;
assign TX_DATA_26_const_net_9              = 4'h0;
assign TX_DATA_27_const_net_9              = 4'h0;
assign TX_DATA_28_const_net_9              = 4'h0;
assign TX_DATA_29_const_net_9              = 4'h0;
assign TX_DATA_30_const_net_9              = 4'h0;
assign TX_DATA_31_const_net_9              = 4'h0;
assign TX_DATA_32_const_net_9              = 4'h0;
assign TX_DATA_33_const_net_9              = 4'h0;
assign TX_DATA_34_const_net_9              = 4'h0;
assign TX_DATA_35_const_net_9              = 4'h0;
assign TX_DATA_36_const_net_9              = 4'h0;
assign TX_DATA_37_const_net_9              = 4'h0;
assign TX_DATA_38_const_net_9              = 4'h0;
assign TX_DATA_39_const_net_9              = 4'h0;
assign TX_DATA_40_const_net_9              = 4'h0;
assign TX_DATA_41_const_net_9              = 4'h0;
assign TX_DATA_42_const_net_9              = 4'h0;
assign TX_DATA_43_const_net_9              = 4'h0;
assign TX_DATA_44_const_net_9              = 4'h0;
assign TX_DATA_45_const_net_9              = 4'h0;
assign TX_DATA_46_const_net_9              = 4'h0;
assign TX_DATA_47_const_net_9              = 4'h0;
assign TX_DATA_48_const_net_9              = 4'h0;
assign TX_DATA_49_const_net_9              = 4'h0;
assign TX_DATA_50_const_net_9              = 4'h0;
assign TX_DATA_51_const_net_9              = 4'h0;
assign TX_DATA_52_const_net_9              = 4'h0;
assign TX_DATA_53_const_net_9              = 4'h0;
assign TX_DATA_54_const_net_9              = 4'h0;
assign TX_DATA_55_const_net_9              = 4'h0;
assign TX_DATA_56_const_net_9              = 4'h0;
assign TX_DATA_57_const_net_9              = 4'h0;
assign TX_DATA_58_const_net_9              = 4'h0;
assign TX_DATA_59_const_net_9              = 4'h0;
assign TX_DATA_60_const_net_9              = 4'h0;
assign TX_DATA_61_const_net_9              = 4'h0;
assign TX_DATA_62_const_net_9              = 4'h0;
assign TX_DATA_63_const_net_9              = 4'h0;
assign TX_DATA_64_const_net_9              = 4'h0;
assign TX_DATA_65_const_net_9              = 4'h0;
assign TX_DATA_66_const_net_9              = 4'h0;
assign TX_DATA_67_const_net_9              = 4'h0;
assign TX_DATA_68_const_net_9              = 4'h0;
assign TX_DATA_69_const_net_9              = 4'h0;
assign TX_DATA_70_const_net_9              = 4'h0;
assign TX_DATA_71_const_net_9              = 4'h0;
assign TX_DATA_72_const_net_9              = 4'h0;
assign TX_DATA_73_const_net_9              = 4'h0;
assign TX_DATA_74_const_net_9              = 4'h0;
assign TX_DATA_75_const_net_9              = 4'h0;
assign TX_DATA_76_const_net_9              = 4'h0;
assign TX_DATA_77_const_net_9              = 4'h0;
assign TX_DATA_78_const_net_9              = 4'h0;
assign TX_DATA_79_const_net_9              = 4'h0;
assign TX_DATA_80_const_net_9              = 4'h0;
assign TX_DATA_81_const_net_9              = 4'h0;
assign TX_DATA_82_const_net_9              = 4'h0;
assign TX_DATA_83_const_net_9              = 4'h0;
assign TX_DATA_84_const_net_9              = 4'h0;
assign TX_DATA_85_const_net_9              = 4'h0;
assign TX_DATA_86_const_net_9              = 4'h0;
assign TX_DATA_87_const_net_9              = 4'h0;
assign TX_DATA_88_const_net_9              = 4'h0;
assign TX_DATA_89_const_net_9              = 4'h0;
assign TX_DATA_90_const_net_9              = 4'h0;
assign TX_DATA_91_const_net_9              = 4'h0;
assign TX_DATA_92_const_net_9              = 4'h0;
assign TX_DATA_93_const_net_9              = 4'h0;
assign TX_DATA_94_const_net_9              = 4'h0;
assign TX_DATA_95_const_net_9              = 4'h0;
assign TX_DATA_96_const_net_9              = 4'h0;
assign TX_DATA_97_const_net_9              = 4'h0;
assign TX_DATA_98_const_net_9              = 4'h0;
assign TX_DATA_99_const_net_9              = 4'h0;
assign TX_DATA_100_const_net_9             = 4'h0;
assign TX_DATA_101_const_net_9             = 4'h0;
assign TX_DATA_102_const_net_9             = 4'h0;
assign TX_DATA_103_const_net_9             = 4'h0;
assign TX_DATA_104_const_net_9             = 4'h0;
assign TX_DATA_105_const_net_9             = 4'h0;
assign TX_DATA_106_const_net_9             = 4'h0;
assign TX_DATA_107_const_net_9             = 4'h0;
assign TX_DATA_108_const_net_9             = 4'h0;
assign TX_DATA_109_const_net_9             = 4'h0;
assign TX_DATA_110_const_net_9             = 4'h0;
assign TX_DATA_111_const_net_9             = 4'h0;
assign TX_DATA_112_const_net_9             = 4'h0;
assign TX_DATA_113_const_net_9             = 4'h0;
assign TX_DATA_114_const_net_9             = 4'h0;
assign TX_DATA_115_const_net_9             = 4'h0;
assign TX_DATA_116_const_net_9             = 4'h0;
assign TX_DATA_117_const_net_9             = 4'h0;
assign TX_DATA_118_const_net_9             = 4'h0;
assign TX_DATA_119_const_net_9             = 4'h0;
assign TX_DATA_120_const_net_9             = 4'h0;
assign TX_DATA_121_const_net_9             = 4'h0;
assign TX_DATA_122_const_net_9             = 4'h0;
assign TX_DATA_123_const_net_9             = 4'h0;
assign TX_DATA_124_const_net_9             = 4'h0;
assign TX_DATA_125_const_net_9             = 4'h0;
assign TX_DATA_126_const_net_9             = 4'h0;
assign TX_DATA_127_const_net_9             = 4'h0;
assign OE_DATA_1_const_net_9               = 4'h0;
assign OE_DATA_2_const_net_9               = 4'h0;
assign OE_DATA_3_const_net_9               = 4'h0;
assign OE_DATA_4_const_net_9               = 4'h0;
assign OE_DATA_5_const_net_9               = 4'h0;
assign OE_DATA_6_const_net_9               = 4'h0;
assign OE_DATA_7_const_net_9               = 4'h0;
assign OE_DATA_8_const_net_9               = 4'h0;
assign OE_DATA_9_const_net_9               = 4'h0;
assign OE_DATA_10_const_net_9              = 4'h0;
assign OE_DATA_11_const_net_9              = 4'h0;
assign OE_DATA_12_const_net_9              = 4'h0;
assign OE_DATA_13_const_net_9              = 4'h0;
assign OE_DATA_14_const_net_9              = 4'h0;
assign OE_DATA_15_const_net_9              = 4'h0;
assign OE_DATA_16_const_net_9              = 4'h0;
assign OE_DATA_17_const_net_9              = 4'h0;
assign OE_DATA_18_const_net_9              = 4'h0;
assign OE_DATA_19_const_net_9              = 4'h0;
assign OE_DATA_20_const_net_9              = 4'h0;
assign OE_DATA_21_const_net_9              = 4'h0;
assign OE_DATA_22_const_net_9              = 4'h0;
assign OE_DATA_23_const_net_9              = 4'h0;
assign OE_DATA_24_const_net_9              = 4'h0;
assign OE_DATA_25_const_net_9              = 4'h0;
assign OE_DATA_26_const_net_9              = 4'h0;
assign OE_DATA_27_const_net_9              = 4'h0;
assign OE_DATA_28_const_net_9              = 4'h0;
assign OE_DATA_29_const_net_9              = 4'h0;
assign OE_DATA_30_const_net_9              = 4'h0;
assign OE_DATA_31_const_net_9              = 4'h0;
assign OE_DATA_32_const_net_9              = 4'h0;
assign OE_DATA_33_const_net_9              = 4'h0;
assign OE_DATA_34_const_net_9              = 4'h0;
assign OE_DATA_35_const_net_9              = 4'h0;
assign OE_DATA_36_const_net_9              = 4'h0;
assign OE_DATA_37_const_net_9              = 4'h0;
assign OE_DATA_38_const_net_9              = 4'h0;
assign OE_DATA_39_const_net_9              = 4'h0;
assign OE_DATA_40_const_net_9              = 4'h0;
assign OE_DATA_41_const_net_9              = 4'h0;
assign OE_DATA_42_const_net_9              = 4'h0;
assign OE_DATA_43_const_net_9              = 4'h0;
assign OE_DATA_44_const_net_9              = 4'h0;
assign OE_DATA_45_const_net_9              = 4'h0;
assign OE_DATA_46_const_net_9              = 4'h0;
assign OE_DATA_47_const_net_9              = 4'h0;
assign OE_DATA_48_const_net_9              = 4'h0;
assign OE_DATA_49_const_net_9              = 4'h0;
assign OE_DATA_50_const_net_9              = 4'h0;
assign OE_DATA_51_const_net_9              = 4'h0;
assign OE_DATA_52_const_net_9              = 4'h0;
assign OE_DATA_53_const_net_9              = 4'h0;
assign OE_DATA_54_const_net_9              = 4'h0;
assign OE_DATA_55_const_net_9              = 4'h0;
assign OE_DATA_56_const_net_9              = 4'h0;
assign OE_DATA_57_const_net_9              = 4'h0;
assign OE_DATA_58_const_net_9              = 4'h0;
assign OE_DATA_59_const_net_9              = 4'h0;
assign OE_DATA_60_const_net_9              = 4'h0;
assign OE_DATA_61_const_net_9              = 4'h0;
assign OE_DATA_62_const_net_9              = 4'h0;
assign OE_DATA_63_const_net_9              = 4'h0;
assign OE_DATA_64_const_net_9              = 4'h0;
assign OE_DATA_65_const_net_9              = 4'h0;
assign OE_DATA_66_const_net_9              = 4'h0;
assign OE_DATA_67_const_net_9              = 4'h0;
assign OE_DATA_68_const_net_9              = 4'h0;
assign OE_DATA_69_const_net_9              = 4'h0;
assign OE_DATA_70_const_net_9              = 4'h0;
assign OE_DATA_71_const_net_9              = 4'h0;
assign OE_DATA_72_const_net_9              = 4'h0;
assign OE_DATA_73_const_net_9              = 4'h0;
assign OE_DATA_74_const_net_9              = 4'h0;
assign OE_DATA_75_const_net_9              = 4'h0;
assign OE_DATA_76_const_net_9              = 4'h0;
assign OE_DATA_77_const_net_9              = 4'h0;
assign OE_DATA_78_const_net_9              = 4'h0;
assign OE_DATA_79_const_net_9              = 4'h0;
assign OE_DATA_80_const_net_9              = 4'h0;
assign OE_DATA_81_const_net_9              = 4'h0;
assign OE_DATA_82_const_net_9              = 4'h0;
assign OE_DATA_83_const_net_9              = 4'h0;
assign OE_DATA_84_const_net_9              = 4'h0;
assign OE_DATA_85_const_net_9              = 4'h0;
assign OE_DATA_86_const_net_9              = 4'h0;
assign OE_DATA_87_const_net_9              = 4'h0;
assign OE_DATA_88_const_net_9              = 4'h0;
assign OE_DATA_89_const_net_9              = 4'h0;
assign OE_DATA_90_const_net_9              = 4'h0;
assign OE_DATA_91_const_net_9              = 4'h0;
assign OE_DATA_92_const_net_9              = 4'h0;
assign OE_DATA_93_const_net_9              = 4'h0;
assign OE_DATA_94_const_net_9              = 4'h0;
assign OE_DATA_95_const_net_9              = 4'h0;
assign OE_DATA_96_const_net_9              = 4'h0;
assign OE_DATA_97_const_net_9              = 4'h0;
assign OE_DATA_98_const_net_9              = 4'h0;
assign OE_DATA_99_const_net_9              = 4'h0;
assign OE_DATA_100_const_net_9             = 4'h0;
assign OE_DATA_101_const_net_9             = 4'h0;
assign OE_DATA_102_const_net_9             = 4'h0;
assign OE_DATA_103_const_net_9             = 4'h0;
assign OE_DATA_104_const_net_9             = 4'h0;
assign OE_DATA_105_const_net_9             = 4'h0;
assign OE_DATA_106_const_net_9             = 4'h0;
assign OE_DATA_107_const_net_9             = 4'h0;
assign OE_DATA_108_const_net_9             = 4'h0;
assign OE_DATA_109_const_net_9             = 4'h0;
assign OE_DATA_110_const_net_9             = 4'h0;
assign OE_DATA_111_const_net_9             = 4'h0;
assign OE_DATA_112_const_net_9             = 4'h0;
assign OE_DATA_113_const_net_9             = 4'h0;
assign OE_DATA_114_const_net_9             = 4'h0;
assign OE_DATA_115_const_net_9             = 4'h0;
assign OE_DATA_116_const_net_9             = 4'h0;
assign OE_DATA_117_const_net_9             = 4'h0;
assign OE_DATA_118_const_net_9             = 4'h0;
assign OE_DATA_119_const_net_9             = 4'h0;
assign OE_DATA_120_const_net_9             = 4'h0;
assign OE_DATA_121_const_net_9             = 4'h0;
assign OE_DATA_122_const_net_9             = 4'h0;
assign OE_DATA_123_const_net_9             = 4'h0;
assign OE_DATA_124_const_net_9             = 4'h0;
assign OE_DATA_125_const_net_9             = 4'h0;
assign OE_DATA_126_const_net_9             = 4'h0;
assign OE_DATA_127_const_net_9             = 4'h0;
assign RX_DQS_90_const_net_10              = 2'h0;
assign FIFO_WR_PTR_const_net_10            = 3'h0;
assign FIFO_RD_PTR_const_net_10            = 3'h0;
assign EYE_MONITOR_LANE_WIDTH_const_net_10 = 3'h0;
assign TX_DATA_1_const_net_7               = 4'h0;
assign TX_DATA_2_const_net_9               = 4'h0;
assign TX_DATA_3_const_net_9               = 4'h0;
assign TX_DATA_4_const_net_9               = 4'h0;
assign TX_DATA_5_const_net_9               = 4'h0;
assign TX_DATA_6_const_net_9               = 4'h0;
assign TX_DATA_7_const_net_9               = 4'h0;
assign TX_DATA_8_const_net_9               = 4'h0;
assign TX_DATA_9_const_net_9               = 4'h0;
assign TX_DATA_10_const_net_9              = 4'h0;
assign TX_DATA_11_const_net_9              = 4'h0;
assign TX_DATA_12_const_net_10             = 4'h0;
assign TX_DATA_13_const_net_10             = 4'h0;
assign TX_DATA_14_const_net_10             = 4'h0;
assign TX_DATA_15_const_net_10             = 4'h0;
assign TX_DATA_16_const_net_10             = 4'h0;
assign TX_DATA_17_const_net_10             = 4'h0;
assign TX_DATA_18_const_net_10             = 4'h0;
assign TX_DATA_19_const_net_10             = 4'h0;
assign TX_DATA_20_const_net_10             = 4'h0;
assign TX_DATA_21_const_net_10             = 4'h0;
assign TX_DATA_22_const_net_10             = 4'h0;
assign TX_DATA_23_const_net_10             = 4'h0;
assign TX_DATA_24_const_net_10             = 4'h0;
assign TX_DATA_25_const_net_10             = 4'h0;
assign TX_DATA_26_const_net_10             = 4'h0;
assign TX_DATA_27_const_net_10             = 4'h0;
assign TX_DATA_28_const_net_10             = 4'h0;
assign TX_DATA_29_const_net_10             = 4'h0;
assign TX_DATA_30_const_net_10             = 4'h0;
assign TX_DATA_31_const_net_10             = 4'h0;
assign TX_DATA_32_const_net_10             = 4'h0;
assign TX_DATA_33_const_net_10             = 4'h0;
assign TX_DATA_34_const_net_10             = 4'h0;
assign TX_DATA_35_const_net_10             = 4'h0;
assign TX_DATA_36_const_net_10             = 4'h0;
assign TX_DATA_37_const_net_10             = 4'h0;
assign TX_DATA_38_const_net_10             = 4'h0;
assign TX_DATA_39_const_net_10             = 4'h0;
assign TX_DATA_40_const_net_10             = 4'h0;
assign TX_DATA_41_const_net_10             = 4'h0;
assign TX_DATA_42_const_net_10             = 4'h0;
assign TX_DATA_43_const_net_10             = 4'h0;
assign TX_DATA_44_const_net_10             = 4'h0;
assign TX_DATA_45_const_net_10             = 4'h0;
assign TX_DATA_46_const_net_10             = 4'h0;
assign TX_DATA_47_const_net_10             = 4'h0;
assign TX_DATA_48_const_net_10             = 4'h0;
assign TX_DATA_49_const_net_10             = 4'h0;
assign TX_DATA_50_const_net_10             = 4'h0;
assign TX_DATA_51_const_net_10             = 4'h0;
assign TX_DATA_52_const_net_10             = 4'h0;
assign TX_DATA_53_const_net_10             = 4'h0;
assign TX_DATA_54_const_net_10             = 4'h0;
assign TX_DATA_55_const_net_10             = 4'h0;
assign TX_DATA_56_const_net_10             = 4'h0;
assign TX_DATA_57_const_net_10             = 4'h0;
assign TX_DATA_58_const_net_10             = 4'h0;
assign TX_DATA_59_const_net_10             = 4'h0;
assign TX_DATA_60_const_net_10             = 4'h0;
assign TX_DATA_61_const_net_10             = 4'h0;
assign TX_DATA_62_const_net_10             = 4'h0;
assign TX_DATA_63_const_net_10             = 4'h0;
assign TX_DATA_64_const_net_10             = 4'h0;
assign TX_DATA_65_const_net_10             = 4'h0;
assign TX_DATA_66_const_net_10             = 4'h0;
assign TX_DATA_67_const_net_10             = 4'h0;
assign TX_DATA_68_const_net_10             = 4'h0;
assign TX_DATA_69_const_net_10             = 4'h0;
assign TX_DATA_70_const_net_10             = 4'h0;
assign TX_DATA_71_const_net_10             = 4'h0;
assign TX_DATA_72_const_net_10             = 4'h0;
assign TX_DATA_73_const_net_10             = 4'h0;
assign TX_DATA_74_const_net_10             = 4'h0;
assign TX_DATA_75_const_net_10             = 4'h0;
assign TX_DATA_76_const_net_10             = 4'h0;
assign TX_DATA_77_const_net_10             = 4'h0;
assign TX_DATA_78_const_net_10             = 4'h0;
assign TX_DATA_79_const_net_10             = 4'h0;
assign TX_DATA_80_const_net_10             = 4'h0;
assign TX_DATA_81_const_net_10             = 4'h0;
assign TX_DATA_82_const_net_10             = 4'h0;
assign TX_DATA_83_const_net_10             = 4'h0;
assign TX_DATA_84_const_net_10             = 4'h0;
assign TX_DATA_85_const_net_10             = 4'h0;
assign TX_DATA_86_const_net_10             = 4'h0;
assign TX_DATA_87_const_net_10             = 4'h0;
assign TX_DATA_88_const_net_10             = 4'h0;
assign TX_DATA_89_const_net_10             = 4'h0;
assign TX_DATA_90_const_net_10             = 4'h0;
assign TX_DATA_91_const_net_10             = 4'h0;
assign TX_DATA_92_const_net_10             = 4'h0;
assign TX_DATA_93_const_net_10             = 4'h0;
assign TX_DATA_94_const_net_10             = 4'h0;
assign TX_DATA_95_const_net_10             = 4'h0;
assign TX_DATA_96_const_net_10             = 4'h0;
assign TX_DATA_97_const_net_10             = 4'h0;
assign TX_DATA_98_const_net_10             = 4'h0;
assign TX_DATA_99_const_net_10             = 4'h0;
assign TX_DATA_100_const_net_10            = 4'h0;
assign TX_DATA_101_const_net_10            = 4'h0;
assign TX_DATA_102_const_net_10            = 4'h0;
assign TX_DATA_103_const_net_10            = 4'h0;
assign TX_DATA_104_const_net_10            = 4'h0;
assign TX_DATA_105_const_net_10            = 4'h0;
assign TX_DATA_106_const_net_10            = 4'h0;
assign TX_DATA_107_const_net_10            = 4'h0;
assign TX_DATA_108_const_net_10            = 4'h0;
assign TX_DATA_109_const_net_10            = 4'h0;
assign TX_DATA_110_const_net_10            = 4'h0;
assign TX_DATA_111_const_net_10            = 4'h0;
assign TX_DATA_112_const_net_10            = 4'h0;
assign TX_DATA_113_const_net_10            = 4'h0;
assign TX_DATA_114_const_net_10            = 4'h0;
assign TX_DATA_115_const_net_10            = 4'h0;
assign TX_DATA_116_const_net_10            = 4'h0;
assign TX_DATA_117_const_net_10            = 4'h0;
assign TX_DATA_118_const_net_10            = 4'h0;
assign TX_DATA_119_const_net_10            = 4'h0;
assign TX_DATA_120_const_net_10            = 4'h0;
assign TX_DATA_121_const_net_10            = 4'h0;
assign TX_DATA_122_const_net_10            = 4'h0;
assign TX_DATA_123_const_net_10            = 4'h0;
assign TX_DATA_124_const_net_10            = 4'h0;
assign TX_DATA_125_const_net_10            = 4'h0;
assign TX_DATA_126_const_net_10            = 4'h0;
assign TX_DATA_127_const_net_10            = 4'h0;
assign OE_DATA_1_const_net_10              = 4'h0;
assign OE_DATA_2_const_net_10              = 4'h0;
assign OE_DATA_3_const_net_10              = 4'h0;
assign OE_DATA_4_const_net_10              = 4'h0;
assign OE_DATA_5_const_net_10              = 4'h0;
assign OE_DATA_6_const_net_10              = 4'h0;
assign OE_DATA_7_const_net_10              = 4'h0;
assign OE_DATA_8_const_net_10              = 4'h0;
assign OE_DATA_9_const_net_10              = 4'h0;
assign OE_DATA_10_const_net_10             = 4'h0;
assign OE_DATA_11_const_net_10             = 4'h0;
assign OE_DATA_12_const_net_10             = 4'h0;
assign OE_DATA_13_const_net_10             = 4'h0;
assign OE_DATA_14_const_net_10             = 4'h0;
assign OE_DATA_15_const_net_10             = 4'h0;
assign OE_DATA_16_const_net_10             = 4'h0;
assign OE_DATA_17_const_net_10             = 4'h0;
assign OE_DATA_18_const_net_10             = 4'h0;
assign OE_DATA_19_const_net_10             = 4'h0;
assign OE_DATA_20_const_net_10             = 4'h0;
assign OE_DATA_21_const_net_10             = 4'h0;
assign OE_DATA_22_const_net_10             = 4'h0;
assign OE_DATA_23_const_net_10             = 4'h0;
assign OE_DATA_24_const_net_10             = 4'h0;
assign OE_DATA_25_const_net_10             = 4'h0;
assign OE_DATA_26_const_net_10             = 4'h0;
assign OE_DATA_27_const_net_10             = 4'h0;
assign OE_DATA_28_const_net_10             = 4'h0;
assign OE_DATA_29_const_net_10             = 4'h0;
assign OE_DATA_30_const_net_10             = 4'h0;
assign OE_DATA_31_const_net_10             = 4'h0;
assign OE_DATA_32_const_net_10             = 4'h0;
assign OE_DATA_33_const_net_10             = 4'h0;
assign OE_DATA_34_const_net_10             = 4'h0;
assign OE_DATA_35_const_net_10             = 4'h0;
assign OE_DATA_36_const_net_10             = 4'h0;
assign OE_DATA_37_const_net_10             = 4'h0;
assign OE_DATA_38_const_net_10             = 4'h0;
assign OE_DATA_39_const_net_10             = 4'h0;
assign OE_DATA_40_const_net_10             = 4'h0;
assign OE_DATA_41_const_net_10             = 4'h0;
assign OE_DATA_42_const_net_10             = 4'h0;
assign OE_DATA_43_const_net_10             = 4'h0;
assign OE_DATA_44_const_net_10             = 4'h0;
assign OE_DATA_45_const_net_10             = 4'h0;
assign OE_DATA_46_const_net_10             = 4'h0;
assign OE_DATA_47_const_net_10             = 4'h0;
assign OE_DATA_48_const_net_10             = 4'h0;
assign OE_DATA_49_const_net_10             = 4'h0;
assign OE_DATA_50_const_net_10             = 4'h0;
assign OE_DATA_51_const_net_10             = 4'h0;
assign OE_DATA_52_const_net_10             = 4'h0;
assign OE_DATA_53_const_net_10             = 4'h0;
assign OE_DATA_54_const_net_10             = 4'h0;
assign OE_DATA_55_const_net_10             = 4'h0;
assign OE_DATA_56_const_net_10             = 4'h0;
assign OE_DATA_57_const_net_10             = 4'h0;
assign OE_DATA_58_const_net_10             = 4'h0;
assign OE_DATA_59_const_net_10             = 4'h0;
assign OE_DATA_60_const_net_10             = 4'h0;
assign OE_DATA_61_const_net_10             = 4'h0;
assign OE_DATA_62_const_net_10             = 4'h0;
assign OE_DATA_63_const_net_10             = 4'h0;
assign OE_DATA_64_const_net_10             = 4'h0;
assign OE_DATA_65_const_net_10             = 4'h0;
assign OE_DATA_66_const_net_10             = 4'h0;
assign OE_DATA_67_const_net_10             = 4'h0;
assign OE_DATA_68_const_net_10             = 4'h0;
assign OE_DATA_69_const_net_10             = 4'h0;
assign OE_DATA_70_const_net_10             = 4'h0;
assign OE_DATA_71_const_net_10             = 4'h0;
assign OE_DATA_72_const_net_10             = 4'h0;
assign OE_DATA_73_const_net_10             = 4'h0;
assign OE_DATA_74_const_net_10             = 4'h0;
assign OE_DATA_75_const_net_10             = 4'h0;
assign OE_DATA_76_const_net_10             = 4'h0;
assign OE_DATA_77_const_net_10             = 4'h0;
assign OE_DATA_78_const_net_10             = 4'h0;
assign OE_DATA_79_const_net_10             = 4'h0;
assign OE_DATA_80_const_net_10             = 4'h0;
assign OE_DATA_81_const_net_10             = 4'h0;
assign OE_DATA_82_const_net_10             = 4'h0;
assign OE_DATA_83_const_net_10             = 4'h0;
assign OE_DATA_84_const_net_10             = 4'h0;
assign OE_DATA_85_const_net_10             = 4'h0;
assign OE_DATA_86_const_net_10             = 4'h0;
assign OE_DATA_87_const_net_10             = 4'h0;
assign OE_DATA_88_const_net_10             = 4'h0;
assign OE_DATA_89_const_net_10             = 4'h0;
assign OE_DATA_90_const_net_10             = 4'h0;
assign OE_DATA_91_const_net_10             = 4'h0;
assign OE_DATA_92_const_net_10             = 4'h0;
assign OE_DATA_93_const_net_10             = 4'h0;
assign OE_DATA_94_const_net_10             = 4'h0;
assign OE_DATA_95_const_net_10             = 4'h0;
assign OE_DATA_96_const_net_10             = 4'h0;
assign OE_DATA_97_const_net_10             = 4'h0;
assign OE_DATA_98_const_net_10             = 4'h0;
assign OE_DATA_99_const_net_10             = 4'h0;
assign OE_DATA_100_const_net_10            = 4'h0;
assign OE_DATA_101_const_net_10            = 4'h0;
assign OE_DATA_102_const_net_10            = 4'h0;
assign OE_DATA_103_const_net_10            = 4'h0;
assign OE_DATA_104_const_net_10            = 4'h0;
assign OE_DATA_105_const_net_10            = 4'h0;
assign OE_DATA_106_const_net_10            = 4'h0;
assign OE_DATA_107_const_net_10            = 4'h0;
assign OE_DATA_108_const_net_10            = 4'h0;
assign OE_DATA_109_const_net_10            = 4'h0;
assign OE_DATA_110_const_net_10            = 4'h0;
assign OE_DATA_111_const_net_10            = 4'h0;
assign OE_DATA_112_const_net_10            = 4'h0;
assign OE_DATA_113_const_net_10            = 4'h0;
assign OE_DATA_114_const_net_10            = 4'h0;
assign OE_DATA_115_const_net_10            = 4'h0;
assign OE_DATA_116_const_net_10            = 4'h0;
assign OE_DATA_117_const_net_10            = 4'h0;
assign OE_DATA_118_const_net_10            = 4'h0;
assign OE_DATA_119_const_net_10            = 4'h0;
assign OE_DATA_120_const_net_10            = 4'h0;
assign OE_DATA_121_const_net_10            = 4'h0;
assign OE_DATA_122_const_net_10            = 4'h0;
assign OE_DATA_123_const_net_10            = 4'h0;
assign OE_DATA_124_const_net_10            = 4'h0;
assign OE_DATA_125_const_net_10            = 4'h0;
assign OE_DATA_126_const_net_10            = 4'h0;
assign OE_DATA_127_const_net_10            = 4'h0;
assign RX_DQS_90_const_net_11              = 2'h0;
assign FIFO_WR_PTR_const_net_11            = 3'h0;
assign FIFO_RD_PTR_const_net_11            = 3'h0;
assign EYE_MONITOR_LANE_WIDTH_const_net_11 = 3'h0;
assign TX_DATA_1_const_net_8               = 4'h0;
assign TX_DATA_2_const_net_10              = 4'h0;
assign TX_DATA_3_const_net_10              = 4'h0;
assign TX_DATA_4_const_net_10              = 4'h0;
assign TX_DATA_5_const_net_10              = 4'h0;
assign TX_DATA_6_const_net_10              = 4'h0;
assign TX_DATA_7_const_net_10              = 4'h0;
assign TX_DATA_8_const_net_10              = 4'h0;
assign TX_DATA_9_const_net_10              = 4'h0;
assign TX_DATA_10_const_net_10             = 4'h0;
assign TX_DATA_11_const_net_10             = 4'h0;
assign TX_DATA_12_const_net_11             = 4'h0;
assign TX_DATA_13_const_net_11             = 4'h0;
assign TX_DATA_14_const_net_11             = 4'h0;
assign TX_DATA_15_const_net_11             = 4'h0;
assign TX_DATA_16_const_net_11             = 4'h0;
assign TX_DATA_17_const_net_11             = 4'h0;
assign TX_DATA_18_const_net_11             = 4'h0;
assign TX_DATA_19_const_net_11             = 4'h0;
assign TX_DATA_20_const_net_11             = 4'h0;
assign TX_DATA_21_const_net_11             = 4'h0;
assign TX_DATA_22_const_net_11             = 4'h0;
assign TX_DATA_23_const_net_11             = 4'h0;
assign TX_DATA_24_const_net_11             = 4'h0;
assign TX_DATA_25_const_net_11             = 4'h0;
assign TX_DATA_26_const_net_11             = 4'h0;
assign TX_DATA_27_const_net_11             = 4'h0;
assign TX_DATA_28_const_net_11             = 4'h0;
assign TX_DATA_29_const_net_11             = 4'h0;
assign TX_DATA_30_const_net_11             = 4'h0;
assign TX_DATA_31_const_net_11             = 4'h0;
assign TX_DATA_32_const_net_11             = 4'h0;
assign TX_DATA_33_const_net_11             = 4'h0;
assign TX_DATA_34_const_net_11             = 4'h0;
assign TX_DATA_35_const_net_11             = 4'h0;
assign TX_DATA_36_const_net_11             = 4'h0;
assign TX_DATA_37_const_net_11             = 4'h0;
assign TX_DATA_38_const_net_11             = 4'h0;
assign TX_DATA_39_const_net_11             = 4'h0;
assign TX_DATA_40_const_net_11             = 4'h0;
assign TX_DATA_41_const_net_11             = 4'h0;
assign TX_DATA_42_const_net_11             = 4'h0;
assign TX_DATA_43_const_net_11             = 4'h0;
assign TX_DATA_44_const_net_11             = 4'h0;
assign TX_DATA_45_const_net_11             = 4'h0;
assign TX_DATA_46_const_net_11             = 4'h0;
assign TX_DATA_47_const_net_11             = 4'h0;
assign TX_DATA_48_const_net_11             = 4'h0;
assign TX_DATA_49_const_net_11             = 4'h0;
assign TX_DATA_50_const_net_11             = 4'h0;
assign TX_DATA_51_const_net_11             = 4'h0;
assign TX_DATA_52_const_net_11             = 4'h0;
assign TX_DATA_53_const_net_11             = 4'h0;
assign TX_DATA_54_const_net_11             = 4'h0;
assign TX_DATA_55_const_net_11             = 4'h0;
assign TX_DATA_56_const_net_11             = 4'h0;
assign TX_DATA_57_const_net_11             = 4'h0;
assign TX_DATA_58_const_net_11             = 4'h0;
assign TX_DATA_59_const_net_11             = 4'h0;
assign TX_DATA_60_const_net_11             = 4'h0;
assign TX_DATA_61_const_net_11             = 4'h0;
assign TX_DATA_62_const_net_11             = 4'h0;
assign TX_DATA_63_const_net_11             = 4'h0;
assign TX_DATA_64_const_net_11             = 4'h0;
assign TX_DATA_65_const_net_11             = 4'h0;
assign TX_DATA_66_const_net_11             = 4'h0;
assign TX_DATA_67_const_net_11             = 4'h0;
assign TX_DATA_68_const_net_11             = 4'h0;
assign TX_DATA_69_const_net_11             = 4'h0;
assign TX_DATA_70_const_net_11             = 4'h0;
assign TX_DATA_71_const_net_11             = 4'h0;
assign TX_DATA_72_const_net_11             = 4'h0;
assign TX_DATA_73_const_net_11             = 4'h0;
assign TX_DATA_74_const_net_11             = 4'h0;
assign TX_DATA_75_const_net_11             = 4'h0;
assign TX_DATA_76_const_net_11             = 4'h0;
assign TX_DATA_77_const_net_11             = 4'h0;
assign TX_DATA_78_const_net_11             = 4'h0;
assign TX_DATA_79_const_net_11             = 4'h0;
assign TX_DATA_80_const_net_11             = 4'h0;
assign TX_DATA_81_const_net_11             = 4'h0;
assign TX_DATA_82_const_net_11             = 4'h0;
assign TX_DATA_83_const_net_11             = 4'h0;
assign TX_DATA_84_const_net_11             = 4'h0;
assign TX_DATA_85_const_net_11             = 4'h0;
assign TX_DATA_86_const_net_11             = 4'h0;
assign TX_DATA_87_const_net_11             = 4'h0;
assign TX_DATA_88_const_net_11             = 4'h0;
assign TX_DATA_89_const_net_11             = 4'h0;
assign TX_DATA_90_const_net_11             = 4'h0;
assign TX_DATA_91_const_net_11             = 4'h0;
assign TX_DATA_92_const_net_11             = 4'h0;
assign TX_DATA_93_const_net_11             = 4'h0;
assign TX_DATA_94_const_net_11             = 4'h0;
assign TX_DATA_95_const_net_11             = 4'h0;
assign TX_DATA_96_const_net_11             = 4'h0;
assign TX_DATA_97_const_net_11             = 4'h0;
assign TX_DATA_98_const_net_11             = 4'h0;
assign TX_DATA_99_const_net_11             = 4'h0;
assign TX_DATA_100_const_net_11            = 4'h0;
assign TX_DATA_101_const_net_11            = 4'h0;
assign TX_DATA_102_const_net_11            = 4'h0;
assign TX_DATA_103_const_net_11            = 4'h0;
assign TX_DATA_104_const_net_11            = 4'h0;
assign TX_DATA_105_const_net_11            = 4'h0;
assign TX_DATA_106_const_net_11            = 4'h0;
assign TX_DATA_107_const_net_11            = 4'h0;
assign TX_DATA_108_const_net_11            = 4'h0;
assign TX_DATA_109_const_net_11            = 4'h0;
assign TX_DATA_110_const_net_11            = 4'h0;
assign TX_DATA_111_const_net_11            = 4'h0;
assign TX_DATA_112_const_net_11            = 4'h0;
assign TX_DATA_113_const_net_11            = 4'h0;
assign TX_DATA_114_const_net_11            = 4'h0;
assign TX_DATA_115_const_net_11            = 4'h0;
assign TX_DATA_116_const_net_11            = 4'h0;
assign TX_DATA_117_const_net_11            = 4'h0;
assign TX_DATA_118_const_net_11            = 4'h0;
assign TX_DATA_119_const_net_11            = 4'h0;
assign TX_DATA_120_const_net_11            = 4'h0;
assign TX_DATA_121_const_net_11            = 4'h0;
assign TX_DATA_122_const_net_11            = 4'h0;
assign TX_DATA_123_const_net_11            = 4'h0;
assign TX_DATA_124_const_net_11            = 4'h0;
assign TX_DATA_125_const_net_11            = 4'h0;
assign TX_DATA_126_const_net_11            = 4'h0;
assign TX_DATA_127_const_net_11            = 4'h0;
assign OE_DATA_1_const_net_11              = 4'h0;
assign OE_DATA_2_const_net_11              = 4'h0;
assign OE_DATA_3_const_net_11              = 4'h0;
assign OE_DATA_4_const_net_11              = 4'h0;
assign OE_DATA_5_const_net_11              = 4'h0;
assign OE_DATA_6_const_net_11              = 4'h0;
assign OE_DATA_7_const_net_11              = 4'h0;
assign OE_DATA_8_const_net_11              = 4'h0;
assign OE_DATA_9_const_net_11              = 4'h0;
assign OE_DATA_10_const_net_11             = 4'h0;
assign OE_DATA_11_const_net_11             = 4'h0;
assign OE_DATA_12_const_net_11             = 4'h0;
assign OE_DATA_13_const_net_11             = 4'h0;
assign OE_DATA_14_const_net_11             = 4'h0;
assign OE_DATA_15_const_net_11             = 4'h0;
assign OE_DATA_16_const_net_11             = 4'h0;
assign OE_DATA_17_const_net_11             = 4'h0;
assign OE_DATA_18_const_net_11             = 4'h0;
assign OE_DATA_19_const_net_11             = 4'h0;
assign OE_DATA_20_const_net_11             = 4'h0;
assign OE_DATA_21_const_net_11             = 4'h0;
assign OE_DATA_22_const_net_11             = 4'h0;
assign OE_DATA_23_const_net_11             = 4'h0;
assign OE_DATA_24_const_net_11             = 4'h0;
assign OE_DATA_25_const_net_11             = 4'h0;
assign OE_DATA_26_const_net_11             = 4'h0;
assign OE_DATA_27_const_net_11             = 4'h0;
assign OE_DATA_28_const_net_11             = 4'h0;
assign OE_DATA_29_const_net_11             = 4'h0;
assign OE_DATA_30_const_net_11             = 4'h0;
assign OE_DATA_31_const_net_11             = 4'h0;
assign OE_DATA_32_const_net_11             = 4'h0;
assign OE_DATA_33_const_net_11             = 4'h0;
assign OE_DATA_34_const_net_11             = 4'h0;
assign OE_DATA_35_const_net_11             = 4'h0;
assign OE_DATA_36_const_net_11             = 4'h0;
assign OE_DATA_37_const_net_11             = 4'h0;
assign OE_DATA_38_const_net_11             = 4'h0;
assign OE_DATA_39_const_net_11             = 4'h0;
assign OE_DATA_40_const_net_11             = 4'h0;
assign OE_DATA_41_const_net_11             = 4'h0;
assign OE_DATA_42_const_net_11             = 4'h0;
assign OE_DATA_43_const_net_11             = 4'h0;
assign OE_DATA_44_const_net_11             = 4'h0;
assign OE_DATA_45_const_net_11             = 4'h0;
assign OE_DATA_46_const_net_11             = 4'h0;
assign OE_DATA_47_const_net_11             = 4'h0;
assign OE_DATA_48_const_net_11             = 4'h0;
assign OE_DATA_49_const_net_11             = 4'h0;
assign OE_DATA_50_const_net_11             = 4'h0;
assign OE_DATA_51_const_net_11             = 4'h0;
assign OE_DATA_52_const_net_11             = 4'h0;
assign OE_DATA_53_const_net_11             = 4'h0;
assign OE_DATA_54_const_net_11             = 4'h0;
assign OE_DATA_55_const_net_11             = 4'h0;
assign OE_DATA_56_const_net_11             = 4'h0;
assign OE_DATA_57_const_net_11             = 4'h0;
assign OE_DATA_58_const_net_11             = 4'h0;
assign OE_DATA_59_const_net_11             = 4'h0;
assign OE_DATA_60_const_net_11             = 4'h0;
assign OE_DATA_61_const_net_11             = 4'h0;
assign OE_DATA_62_const_net_11             = 4'h0;
assign OE_DATA_63_const_net_11             = 4'h0;
assign OE_DATA_64_const_net_11             = 4'h0;
assign OE_DATA_65_const_net_11             = 4'h0;
assign OE_DATA_66_const_net_11             = 4'h0;
assign OE_DATA_67_const_net_11             = 4'h0;
assign OE_DATA_68_const_net_11             = 4'h0;
assign OE_DATA_69_const_net_11             = 4'h0;
assign OE_DATA_70_const_net_11             = 4'h0;
assign OE_DATA_71_const_net_11             = 4'h0;
assign OE_DATA_72_const_net_11             = 4'h0;
assign OE_DATA_73_const_net_11             = 4'h0;
assign OE_DATA_74_const_net_11             = 4'h0;
assign OE_DATA_75_const_net_11             = 4'h0;
assign OE_DATA_76_const_net_11             = 4'h0;
assign OE_DATA_77_const_net_11             = 4'h0;
assign OE_DATA_78_const_net_11             = 4'h0;
assign OE_DATA_79_const_net_11             = 4'h0;
assign OE_DATA_80_const_net_11             = 4'h0;
assign OE_DATA_81_const_net_11             = 4'h0;
assign OE_DATA_82_const_net_11             = 4'h0;
assign OE_DATA_83_const_net_11             = 4'h0;
assign OE_DATA_84_const_net_11             = 4'h0;
assign OE_DATA_85_const_net_11             = 4'h0;
assign OE_DATA_86_const_net_11             = 4'h0;
assign OE_DATA_87_const_net_11             = 4'h0;
assign OE_DATA_88_const_net_11             = 4'h0;
assign OE_DATA_89_const_net_11             = 4'h0;
assign OE_DATA_90_const_net_11             = 4'h0;
assign OE_DATA_91_const_net_11             = 4'h0;
assign OE_DATA_92_const_net_11             = 4'h0;
assign OE_DATA_93_const_net_11             = 4'h0;
assign OE_DATA_94_const_net_11             = 4'h0;
assign OE_DATA_95_const_net_11             = 4'h0;
assign OE_DATA_96_const_net_11             = 4'h0;
assign OE_DATA_97_const_net_11             = 4'h0;
assign OE_DATA_98_const_net_11             = 4'h0;
assign OE_DATA_99_const_net_11             = 4'h0;
assign OE_DATA_100_const_net_11            = 4'h0;
assign OE_DATA_101_const_net_11            = 4'h0;
assign OE_DATA_102_const_net_11            = 4'h0;
assign OE_DATA_103_const_net_11            = 4'h0;
assign OE_DATA_104_const_net_11            = 4'h0;
assign OE_DATA_105_const_net_11            = 4'h0;
assign OE_DATA_106_const_net_11            = 4'h0;
assign OE_DATA_107_const_net_11            = 4'h0;
assign OE_DATA_108_const_net_11            = 4'h0;
assign OE_DATA_109_const_net_11            = 4'h0;
assign OE_DATA_110_const_net_11            = 4'h0;
assign OE_DATA_111_const_net_11            = 4'h0;
assign OE_DATA_112_const_net_11            = 4'h0;
assign OE_DATA_113_const_net_11            = 4'h0;
assign OE_DATA_114_const_net_11            = 4'h0;
assign OE_DATA_115_const_net_11            = 4'h0;
assign OE_DATA_116_const_net_11            = 4'h0;
assign OE_DATA_117_const_net_11            = 4'h0;
assign OE_DATA_118_const_net_11            = 4'h0;
assign OE_DATA_119_const_net_11            = 4'h0;
assign OE_DATA_120_const_net_11            = 4'h0;
assign OE_DATA_121_const_net_11            = 4'h0;
assign OE_DATA_122_const_net_11            = 4'h0;
assign OE_DATA_123_const_net_11            = 4'h0;
assign OE_DATA_124_const_net_11            = 4'h0;
assign OE_DATA_125_const_net_11            = 4'h0;
assign OE_DATA_126_const_net_11            = 4'h0;
assign OE_DATA_127_const_net_11            = 4'h0;
assign RX_DQS_90_const_net_12              = 2'h0;
assign FIFO_WR_PTR_const_net_12            = 3'h0;
assign FIFO_RD_PTR_const_net_12            = 3'h0;
assign EYE_MONITOR_LANE_WIDTH_const_net_12 = 3'h0;
assign TX_DATA_0_const_net_9               = 8'h00;
assign TX_DATA_1_const_net_9               = 8'h00;
assign TX_DATA_2_const_net_11              = 8'h00;
assign TX_DATA_3_const_net_11              = 8'h00;
assign TX_DATA_4_const_net_11              = 8'h00;
assign TX_DATA_5_const_net_11              = 8'h00;
assign TX_DATA_6_const_net_11              = 8'h00;
assign TX_DATA_7_const_net_11              = 8'h00;
assign TX_DATA_8_const_net_11              = 8'h00;
assign TX_DATA_9_const_net_11              = 8'h00;
assign TX_DATA_10_const_net_11             = 8'h00;
assign TX_DATA_11_const_net_11             = 8'h00;
assign TX_DATA_12_const_net_12             = 8'h00;
assign TX_DATA_13_const_net_12             = 8'h00;
assign TX_DATA_14_const_net_12             = 8'h00;
assign TX_DATA_15_const_net_12             = 8'h00;
assign TX_DATA_16_const_net_12             = 8'h00;
assign TX_DATA_17_const_net_12             = 8'h00;
assign TX_DATA_18_const_net_12             = 8'h00;
assign TX_DATA_19_const_net_12             = 8'h00;
assign TX_DATA_20_const_net_12             = 8'h00;
assign TX_DATA_21_const_net_12             = 8'h00;
assign TX_DATA_22_const_net_12             = 8'h00;
assign TX_DATA_23_const_net_12             = 8'h00;
assign TX_DATA_24_const_net_12             = 8'h00;
assign TX_DATA_25_const_net_12             = 8'h00;
assign TX_DATA_26_const_net_12             = 8'h00;
assign TX_DATA_27_const_net_12             = 8'h00;
assign TX_DATA_28_const_net_12             = 8'h00;
assign TX_DATA_29_const_net_12             = 8'h00;
assign TX_DATA_30_const_net_12             = 8'h00;
assign TX_DATA_31_const_net_12             = 8'h00;
assign TX_DATA_32_const_net_12             = 8'h00;
assign TX_DATA_33_const_net_12             = 8'h00;
assign TX_DATA_34_const_net_12             = 8'h00;
assign TX_DATA_35_const_net_12             = 8'h00;
assign TX_DATA_36_const_net_12             = 8'h00;
assign TX_DATA_37_const_net_12             = 8'h00;
assign TX_DATA_38_const_net_12             = 8'h00;
assign TX_DATA_39_const_net_12             = 8'h00;
assign TX_DATA_40_const_net_12             = 8'h00;
assign TX_DATA_41_const_net_12             = 8'h00;
assign TX_DATA_42_const_net_12             = 8'h00;
assign TX_DATA_43_const_net_12             = 8'h00;
assign TX_DATA_44_const_net_12             = 8'h00;
assign TX_DATA_45_const_net_12             = 8'h00;
assign TX_DATA_46_const_net_12             = 8'h00;
assign TX_DATA_47_const_net_12             = 8'h00;
assign TX_DATA_48_const_net_12             = 8'h00;
assign TX_DATA_49_const_net_12             = 8'h00;
assign TX_DATA_50_const_net_12             = 8'h00;
assign TX_DATA_51_const_net_12             = 8'h00;
assign TX_DATA_52_const_net_12             = 8'h00;
assign TX_DATA_53_const_net_12             = 8'h00;
assign TX_DATA_54_const_net_12             = 8'h00;
assign TX_DATA_55_const_net_12             = 8'h00;
assign TX_DATA_56_const_net_12             = 8'h00;
assign TX_DATA_57_const_net_12             = 8'h00;
assign TX_DATA_58_const_net_12             = 8'h00;
assign TX_DATA_59_const_net_12             = 8'h00;
assign TX_DATA_60_const_net_12             = 8'h00;
assign TX_DATA_61_const_net_12             = 8'h00;
assign TX_DATA_62_const_net_12             = 8'h00;
assign TX_DATA_63_const_net_12             = 8'h00;
assign TX_DATA_64_const_net_12             = 8'h00;
assign TX_DATA_65_const_net_12             = 8'h00;
assign TX_DATA_66_const_net_12             = 8'h00;
assign TX_DATA_67_const_net_12             = 8'h00;
assign TX_DATA_68_const_net_12             = 8'h00;
assign TX_DATA_69_const_net_12             = 8'h00;
assign TX_DATA_70_const_net_12             = 8'h00;
assign TX_DATA_71_const_net_12             = 8'h00;
assign TX_DATA_72_const_net_12             = 8'h00;
assign TX_DATA_73_const_net_12             = 8'h00;
assign TX_DATA_74_const_net_12             = 8'h00;
assign TX_DATA_75_const_net_12             = 8'h00;
assign TX_DATA_76_const_net_12             = 8'h00;
assign TX_DATA_77_const_net_12             = 8'h00;
assign TX_DATA_78_const_net_12             = 8'h00;
assign TX_DATA_79_const_net_12             = 8'h00;
assign TX_DATA_80_const_net_12             = 8'h00;
assign TX_DATA_81_const_net_12             = 8'h00;
assign TX_DATA_82_const_net_12             = 8'h00;
assign TX_DATA_83_const_net_12             = 8'h00;
assign TX_DATA_84_const_net_12             = 8'h00;
assign TX_DATA_85_const_net_12             = 8'h00;
assign TX_DATA_86_const_net_12             = 8'h00;
assign TX_DATA_87_const_net_12             = 8'h00;
assign TX_DATA_88_const_net_12             = 8'h00;
assign TX_DATA_89_const_net_12             = 8'h00;
assign TX_DATA_90_const_net_12             = 8'h00;
assign TX_DATA_91_const_net_12             = 8'h00;
assign TX_DATA_92_const_net_12             = 8'h00;
assign TX_DATA_93_const_net_12             = 8'h00;
assign TX_DATA_94_const_net_12             = 8'h00;
assign TX_DATA_95_const_net_12             = 8'h00;
assign TX_DATA_96_const_net_12             = 8'h00;
assign TX_DATA_97_const_net_12             = 8'h00;
assign TX_DATA_98_const_net_12             = 8'h00;
assign TX_DATA_99_const_net_12             = 8'h00;
assign TX_DATA_100_const_net_12            = 8'h00;
assign TX_DATA_101_const_net_12            = 8'h00;
assign TX_DATA_102_const_net_12            = 8'h00;
assign TX_DATA_103_const_net_12            = 8'h00;
assign TX_DATA_104_const_net_12            = 8'h00;
assign TX_DATA_105_const_net_12            = 8'h00;
assign TX_DATA_106_const_net_12            = 8'h00;
assign TX_DATA_107_const_net_12            = 8'h00;
assign TX_DATA_108_const_net_12            = 8'h00;
assign TX_DATA_109_const_net_12            = 8'h00;
assign TX_DATA_110_const_net_12            = 8'h00;
assign TX_DATA_111_const_net_12            = 8'h00;
assign TX_DATA_112_const_net_12            = 8'h00;
assign TX_DATA_113_const_net_12            = 8'h00;
assign TX_DATA_114_const_net_12            = 8'h00;
assign TX_DATA_115_const_net_12            = 8'h00;
assign TX_DATA_116_const_net_12            = 8'h00;
assign TX_DATA_117_const_net_12            = 8'h00;
assign TX_DATA_118_const_net_12            = 8'h00;
assign TX_DATA_119_const_net_12            = 8'h00;
assign TX_DATA_120_const_net_12            = 8'h00;
assign TX_DATA_121_const_net_12            = 8'h00;
assign TX_DATA_122_const_net_12            = 8'h00;
assign TX_DATA_123_const_net_12            = 8'h00;
assign TX_DATA_124_const_net_12            = 8'h00;
assign TX_DATA_125_const_net_12            = 8'h00;
assign TX_DATA_126_const_net_12            = 8'h00;
assign TX_DATA_127_const_net_12            = 8'h00;
assign OE_DATA_0_const_net_17              = 4'h0;
assign OE_DATA_1_const_net_12              = 4'h0;
assign OE_DATA_2_const_net_12              = 4'h0;
assign OE_DATA_3_const_net_12              = 4'h0;
assign OE_DATA_4_const_net_12              = 4'h0;
assign OE_DATA_5_const_net_12              = 4'h0;
assign OE_DATA_6_const_net_12              = 4'h0;
assign OE_DATA_7_const_net_12              = 4'h0;
assign OE_DATA_8_const_net_12              = 4'h0;
assign OE_DATA_9_const_net_12              = 4'h0;
assign OE_DATA_10_const_net_12             = 4'h0;
assign OE_DATA_11_const_net_12             = 4'h0;
assign OE_DATA_12_const_net_12             = 4'h0;
assign OE_DATA_13_const_net_12             = 4'h0;
assign OE_DATA_14_const_net_12             = 4'h0;
assign OE_DATA_15_const_net_12             = 4'h0;
assign OE_DATA_16_const_net_12             = 4'h0;
assign OE_DATA_17_const_net_12             = 4'h0;
assign OE_DATA_18_const_net_12             = 4'h0;
assign OE_DATA_19_const_net_12             = 4'h0;
assign OE_DATA_20_const_net_12             = 4'h0;
assign OE_DATA_21_const_net_12             = 4'h0;
assign OE_DATA_22_const_net_12             = 4'h0;
assign OE_DATA_23_const_net_12             = 4'h0;
assign OE_DATA_24_const_net_12             = 4'h0;
assign OE_DATA_25_const_net_12             = 4'h0;
assign OE_DATA_26_const_net_12             = 4'h0;
assign OE_DATA_27_const_net_12             = 4'h0;
assign OE_DATA_28_const_net_12             = 4'h0;
assign OE_DATA_29_const_net_12             = 4'h0;
assign OE_DATA_30_const_net_12             = 4'h0;
assign OE_DATA_31_const_net_12             = 4'h0;
assign OE_DATA_32_const_net_12             = 4'h0;
assign OE_DATA_33_const_net_12             = 4'h0;
assign OE_DATA_34_const_net_12             = 4'h0;
assign OE_DATA_35_const_net_12             = 4'h0;
assign OE_DATA_36_const_net_12             = 4'h0;
assign OE_DATA_37_const_net_12             = 4'h0;
assign OE_DATA_38_const_net_12             = 4'h0;
assign OE_DATA_39_const_net_12             = 4'h0;
assign OE_DATA_40_const_net_12             = 4'h0;
assign OE_DATA_41_const_net_12             = 4'h0;
assign OE_DATA_42_const_net_12             = 4'h0;
assign OE_DATA_43_const_net_12             = 4'h0;
assign OE_DATA_44_const_net_12             = 4'h0;
assign OE_DATA_45_const_net_12             = 4'h0;
assign OE_DATA_46_const_net_12             = 4'h0;
assign OE_DATA_47_const_net_12             = 4'h0;
assign OE_DATA_48_const_net_12             = 4'h0;
assign OE_DATA_49_const_net_12             = 4'h0;
assign OE_DATA_50_const_net_12             = 4'h0;
assign OE_DATA_51_const_net_12             = 4'h0;
assign OE_DATA_52_const_net_12             = 4'h0;
assign OE_DATA_53_const_net_12             = 4'h0;
assign OE_DATA_54_const_net_12             = 4'h0;
assign OE_DATA_55_const_net_12             = 4'h0;
assign OE_DATA_56_const_net_12             = 4'h0;
assign OE_DATA_57_const_net_12             = 4'h0;
assign OE_DATA_58_const_net_12             = 4'h0;
assign OE_DATA_59_const_net_12             = 4'h0;
assign OE_DATA_60_const_net_12             = 4'h0;
assign OE_DATA_61_const_net_12             = 4'h0;
assign OE_DATA_62_const_net_12             = 4'h0;
assign OE_DATA_63_const_net_12             = 4'h0;
assign OE_DATA_64_const_net_12             = 4'h0;
assign OE_DATA_65_const_net_12             = 4'h0;
assign OE_DATA_66_const_net_12             = 4'h0;
assign OE_DATA_67_const_net_12             = 4'h0;
assign OE_DATA_68_const_net_12             = 4'h0;
assign OE_DATA_69_const_net_12             = 4'h0;
assign OE_DATA_70_const_net_12             = 4'h0;
assign OE_DATA_71_const_net_12             = 4'h0;
assign OE_DATA_72_const_net_12             = 4'h0;
assign OE_DATA_73_const_net_12             = 4'h0;
assign OE_DATA_74_const_net_12             = 4'h0;
assign OE_DATA_75_const_net_12             = 4'h0;
assign OE_DATA_76_const_net_12             = 4'h0;
assign OE_DATA_77_const_net_12             = 4'h0;
assign OE_DATA_78_const_net_12             = 4'h0;
assign OE_DATA_79_const_net_12             = 4'h0;
assign OE_DATA_80_const_net_12             = 4'h0;
assign OE_DATA_81_const_net_12             = 4'h0;
assign OE_DATA_82_const_net_12             = 4'h0;
assign OE_DATA_83_const_net_12             = 4'h0;
assign OE_DATA_84_const_net_12             = 4'h0;
assign OE_DATA_85_const_net_12             = 4'h0;
assign OE_DATA_86_const_net_12             = 4'h0;
assign OE_DATA_87_const_net_12             = 4'h0;
assign OE_DATA_88_const_net_12             = 4'h0;
assign OE_DATA_89_const_net_12             = 4'h0;
assign OE_DATA_90_const_net_12             = 4'h0;
assign OE_DATA_91_const_net_12             = 4'h0;
assign OE_DATA_92_const_net_12             = 4'h0;
assign OE_DATA_93_const_net_12             = 4'h0;
assign OE_DATA_94_const_net_12             = 4'h0;
assign OE_DATA_95_const_net_12             = 4'h0;
assign OE_DATA_96_const_net_12             = 4'h0;
assign OE_DATA_97_const_net_12             = 4'h0;
assign OE_DATA_98_const_net_12             = 4'h0;
assign OE_DATA_99_const_net_12             = 4'h0;
assign OE_DATA_100_const_net_12            = 4'h0;
assign OE_DATA_101_const_net_12            = 4'h0;
assign OE_DATA_102_const_net_12            = 4'h0;
assign OE_DATA_103_const_net_12            = 4'h0;
assign OE_DATA_104_const_net_12            = 4'h0;
assign OE_DATA_105_const_net_12            = 4'h0;
assign OE_DATA_106_const_net_12            = 4'h0;
assign OE_DATA_107_const_net_12            = 4'h0;
assign OE_DATA_108_const_net_12            = 4'h0;
assign OE_DATA_109_const_net_12            = 4'h0;
assign OE_DATA_110_const_net_12            = 4'h0;
assign OE_DATA_111_const_net_12            = 4'h0;
assign OE_DATA_112_const_net_12            = 4'h0;
assign OE_DATA_113_const_net_12            = 4'h0;
assign OE_DATA_114_const_net_12            = 4'h0;
assign OE_DATA_115_const_net_12            = 4'h0;
assign OE_DATA_116_const_net_12            = 4'h0;
assign OE_DATA_117_const_net_12            = 4'h0;
assign OE_DATA_118_const_net_12            = 4'h0;
assign OE_DATA_119_const_net_12            = 4'h0;
assign OE_DATA_120_const_net_12            = 4'h0;
assign OE_DATA_121_const_net_12            = 4'h0;
assign OE_DATA_122_const_net_12            = 4'h0;
assign OE_DATA_123_const_net_12            = 4'h0;
assign OE_DATA_124_const_net_12            = 4'h0;
assign OE_DATA_125_const_net_12            = 4'h0;
assign OE_DATA_126_const_net_12            = 4'h0;
assign OE_DATA_127_const_net_12            = 4'h0;
assign RX_DQS_90_const_net_13              = 2'h0;
assign FIFO_WR_PTR_const_net_13            = 3'h0;
assign FIFO_RD_PTR_const_net_13            = 3'h0;
assign EYE_MONITOR_LANE_WIDTH_const_net_13 = 3'h0;
assign TX_DATA_1_const_net_10              = 4'h0;
assign TX_DATA_2_const_net_12              = 4'h0;
assign TX_DATA_3_const_net_12              = 4'h0;
assign TX_DATA_4_const_net_12              = 4'h0;
assign TX_DATA_5_const_net_12              = 4'h0;
assign TX_DATA_6_const_net_12              = 4'h0;
assign TX_DATA_7_const_net_12              = 4'h0;
assign TX_DATA_8_const_net_12              = 4'h0;
assign TX_DATA_9_const_net_12              = 4'h0;
assign TX_DATA_10_const_net_12             = 4'h0;
assign TX_DATA_11_const_net_12             = 4'h0;
assign TX_DATA_12_const_net_13             = 4'h0;
assign TX_DATA_13_const_net_13             = 4'h0;
assign TX_DATA_14_const_net_13             = 4'h0;
assign TX_DATA_15_const_net_13             = 4'h0;
assign TX_DATA_16_const_net_13             = 4'h0;
assign TX_DATA_17_const_net_13             = 4'h0;
assign TX_DATA_18_const_net_13             = 4'h0;
assign TX_DATA_19_const_net_13             = 4'h0;
assign TX_DATA_20_const_net_13             = 4'h0;
assign TX_DATA_21_const_net_13             = 4'h0;
assign TX_DATA_22_const_net_13             = 4'h0;
assign TX_DATA_23_const_net_13             = 4'h0;
assign TX_DATA_24_const_net_13             = 4'h0;
assign TX_DATA_25_const_net_13             = 4'h0;
assign TX_DATA_26_const_net_13             = 4'h0;
assign TX_DATA_27_const_net_13             = 4'h0;
assign TX_DATA_28_const_net_13             = 4'h0;
assign TX_DATA_29_const_net_13             = 4'h0;
assign TX_DATA_30_const_net_13             = 4'h0;
assign TX_DATA_31_const_net_13             = 4'h0;
assign TX_DATA_32_const_net_13             = 4'h0;
assign TX_DATA_33_const_net_13             = 4'h0;
assign TX_DATA_34_const_net_13             = 4'h0;
assign TX_DATA_35_const_net_13             = 4'h0;
assign TX_DATA_36_const_net_13             = 4'h0;
assign TX_DATA_37_const_net_13             = 4'h0;
assign TX_DATA_38_const_net_13             = 4'h0;
assign TX_DATA_39_const_net_13             = 4'h0;
assign TX_DATA_40_const_net_13             = 4'h0;
assign TX_DATA_41_const_net_13             = 4'h0;
assign TX_DATA_42_const_net_13             = 4'h0;
assign TX_DATA_43_const_net_13             = 4'h0;
assign TX_DATA_44_const_net_13             = 4'h0;
assign TX_DATA_45_const_net_13             = 4'h0;
assign TX_DATA_46_const_net_13             = 4'h0;
assign TX_DATA_47_const_net_13             = 4'h0;
assign TX_DATA_48_const_net_13             = 4'h0;
assign TX_DATA_49_const_net_13             = 4'h0;
assign TX_DATA_50_const_net_13             = 4'h0;
assign TX_DATA_51_const_net_13             = 4'h0;
assign TX_DATA_52_const_net_13             = 4'h0;
assign TX_DATA_53_const_net_13             = 4'h0;
assign TX_DATA_54_const_net_13             = 4'h0;
assign TX_DATA_55_const_net_13             = 4'h0;
assign TX_DATA_56_const_net_13             = 4'h0;
assign TX_DATA_57_const_net_13             = 4'h0;
assign TX_DATA_58_const_net_13             = 4'h0;
assign TX_DATA_59_const_net_13             = 4'h0;
assign TX_DATA_60_const_net_13             = 4'h0;
assign TX_DATA_61_const_net_13             = 4'h0;
assign TX_DATA_62_const_net_13             = 4'h0;
assign TX_DATA_63_const_net_13             = 4'h0;
assign TX_DATA_64_const_net_13             = 4'h0;
assign TX_DATA_65_const_net_13             = 4'h0;
assign TX_DATA_66_const_net_13             = 4'h0;
assign TX_DATA_67_const_net_13             = 4'h0;
assign TX_DATA_68_const_net_13             = 4'h0;
assign TX_DATA_69_const_net_13             = 4'h0;
assign TX_DATA_70_const_net_13             = 4'h0;
assign TX_DATA_71_const_net_13             = 4'h0;
assign TX_DATA_72_const_net_13             = 4'h0;
assign TX_DATA_73_const_net_13             = 4'h0;
assign TX_DATA_74_const_net_13             = 4'h0;
assign TX_DATA_75_const_net_13             = 4'h0;
assign TX_DATA_76_const_net_13             = 4'h0;
assign TX_DATA_77_const_net_13             = 4'h0;
assign TX_DATA_78_const_net_13             = 4'h0;
assign TX_DATA_79_const_net_13             = 4'h0;
assign TX_DATA_80_const_net_13             = 4'h0;
assign TX_DATA_81_const_net_13             = 4'h0;
assign TX_DATA_82_const_net_13             = 4'h0;
assign TX_DATA_83_const_net_13             = 4'h0;
assign TX_DATA_84_const_net_13             = 4'h0;
assign TX_DATA_85_const_net_13             = 4'h0;
assign TX_DATA_86_const_net_13             = 4'h0;
assign TX_DATA_87_const_net_13             = 4'h0;
assign TX_DATA_88_const_net_13             = 4'h0;
assign TX_DATA_89_const_net_13             = 4'h0;
assign TX_DATA_90_const_net_13             = 4'h0;
assign TX_DATA_91_const_net_13             = 4'h0;
assign TX_DATA_92_const_net_13             = 4'h0;
assign TX_DATA_93_const_net_13             = 4'h0;
assign TX_DATA_94_const_net_13             = 4'h0;
assign TX_DATA_95_const_net_13             = 4'h0;
assign TX_DATA_96_const_net_13             = 4'h0;
assign TX_DATA_97_const_net_13             = 4'h0;
assign TX_DATA_98_const_net_13             = 4'h0;
assign TX_DATA_99_const_net_13             = 4'h0;
assign TX_DATA_100_const_net_13            = 4'h0;
assign TX_DATA_101_const_net_13            = 4'h0;
assign TX_DATA_102_const_net_13            = 4'h0;
assign TX_DATA_103_const_net_13            = 4'h0;
assign TX_DATA_104_const_net_13            = 4'h0;
assign TX_DATA_105_const_net_13            = 4'h0;
assign TX_DATA_106_const_net_13            = 4'h0;
assign TX_DATA_107_const_net_13            = 4'h0;
assign TX_DATA_108_const_net_13            = 4'h0;
assign TX_DATA_109_const_net_13            = 4'h0;
assign TX_DATA_110_const_net_13            = 4'h0;
assign TX_DATA_111_const_net_13            = 4'h0;
assign TX_DATA_112_const_net_13            = 4'h0;
assign TX_DATA_113_const_net_13            = 4'h0;
assign TX_DATA_114_const_net_13            = 4'h0;
assign TX_DATA_115_const_net_13            = 4'h0;
assign TX_DATA_116_const_net_13            = 4'h0;
assign TX_DATA_117_const_net_13            = 4'h0;
assign TX_DATA_118_const_net_13            = 4'h0;
assign TX_DATA_119_const_net_13            = 4'h0;
assign TX_DATA_120_const_net_13            = 4'h0;
assign TX_DATA_121_const_net_13            = 4'h0;
assign TX_DATA_122_const_net_13            = 4'h0;
assign TX_DATA_123_const_net_13            = 4'h0;
assign TX_DATA_124_const_net_13            = 4'h0;
assign TX_DATA_125_const_net_13            = 4'h0;
assign TX_DATA_126_const_net_13            = 4'h0;
assign TX_DATA_127_const_net_13            = 4'h0;
assign OE_DATA_1_const_net_13              = 4'h0;
assign OE_DATA_2_const_net_13              = 4'h0;
assign OE_DATA_3_const_net_13              = 4'h0;
assign OE_DATA_4_const_net_13              = 4'h0;
assign OE_DATA_5_const_net_13              = 4'h0;
assign OE_DATA_6_const_net_13              = 4'h0;
assign OE_DATA_7_const_net_13              = 4'h0;
assign OE_DATA_8_const_net_13              = 4'h0;
assign OE_DATA_9_const_net_13              = 4'h0;
assign OE_DATA_10_const_net_13             = 4'h0;
assign OE_DATA_11_const_net_13             = 4'h0;
assign OE_DATA_12_const_net_13             = 4'h0;
assign OE_DATA_13_const_net_13             = 4'h0;
assign OE_DATA_14_const_net_13             = 4'h0;
assign OE_DATA_15_const_net_13             = 4'h0;
assign OE_DATA_16_const_net_13             = 4'h0;
assign OE_DATA_17_const_net_13             = 4'h0;
assign OE_DATA_18_const_net_13             = 4'h0;
assign OE_DATA_19_const_net_13             = 4'h0;
assign OE_DATA_20_const_net_13             = 4'h0;
assign OE_DATA_21_const_net_13             = 4'h0;
assign OE_DATA_22_const_net_13             = 4'h0;
assign OE_DATA_23_const_net_13             = 4'h0;
assign OE_DATA_24_const_net_13             = 4'h0;
assign OE_DATA_25_const_net_13             = 4'h0;
assign OE_DATA_26_const_net_13             = 4'h0;
assign OE_DATA_27_const_net_13             = 4'h0;
assign OE_DATA_28_const_net_13             = 4'h0;
assign OE_DATA_29_const_net_13             = 4'h0;
assign OE_DATA_30_const_net_13             = 4'h0;
assign OE_DATA_31_const_net_13             = 4'h0;
assign OE_DATA_32_const_net_13             = 4'h0;
assign OE_DATA_33_const_net_13             = 4'h0;
assign OE_DATA_34_const_net_13             = 4'h0;
assign OE_DATA_35_const_net_13             = 4'h0;
assign OE_DATA_36_const_net_13             = 4'h0;
assign OE_DATA_37_const_net_13             = 4'h0;
assign OE_DATA_38_const_net_13             = 4'h0;
assign OE_DATA_39_const_net_13             = 4'h0;
assign OE_DATA_40_const_net_13             = 4'h0;
assign OE_DATA_41_const_net_13             = 4'h0;
assign OE_DATA_42_const_net_13             = 4'h0;
assign OE_DATA_43_const_net_13             = 4'h0;
assign OE_DATA_44_const_net_13             = 4'h0;
assign OE_DATA_45_const_net_13             = 4'h0;
assign OE_DATA_46_const_net_13             = 4'h0;
assign OE_DATA_47_const_net_13             = 4'h0;
assign OE_DATA_48_const_net_13             = 4'h0;
assign OE_DATA_49_const_net_13             = 4'h0;
assign OE_DATA_50_const_net_13             = 4'h0;
assign OE_DATA_51_const_net_13             = 4'h0;
assign OE_DATA_52_const_net_13             = 4'h0;
assign OE_DATA_53_const_net_13             = 4'h0;
assign OE_DATA_54_const_net_13             = 4'h0;
assign OE_DATA_55_const_net_13             = 4'h0;
assign OE_DATA_56_const_net_13             = 4'h0;
assign OE_DATA_57_const_net_13             = 4'h0;
assign OE_DATA_58_const_net_13             = 4'h0;
assign OE_DATA_59_const_net_13             = 4'h0;
assign OE_DATA_60_const_net_13             = 4'h0;
assign OE_DATA_61_const_net_13             = 4'h0;
assign OE_DATA_62_const_net_13             = 4'h0;
assign OE_DATA_63_const_net_13             = 4'h0;
assign OE_DATA_64_const_net_13             = 4'h0;
assign OE_DATA_65_const_net_13             = 4'h0;
assign OE_DATA_66_const_net_13             = 4'h0;
assign OE_DATA_67_const_net_13             = 4'h0;
assign OE_DATA_68_const_net_13             = 4'h0;
assign OE_DATA_69_const_net_13             = 4'h0;
assign OE_DATA_70_const_net_13             = 4'h0;
assign OE_DATA_71_const_net_13             = 4'h0;
assign OE_DATA_72_const_net_13             = 4'h0;
assign OE_DATA_73_const_net_13             = 4'h0;
assign OE_DATA_74_const_net_13             = 4'h0;
assign OE_DATA_75_const_net_13             = 4'h0;
assign OE_DATA_76_const_net_13             = 4'h0;
assign OE_DATA_77_const_net_13             = 4'h0;
assign OE_DATA_78_const_net_13             = 4'h0;
assign OE_DATA_79_const_net_13             = 4'h0;
assign OE_DATA_80_const_net_13             = 4'h0;
assign OE_DATA_81_const_net_13             = 4'h0;
assign OE_DATA_82_const_net_13             = 4'h0;
assign OE_DATA_83_const_net_13             = 4'h0;
assign OE_DATA_84_const_net_13             = 4'h0;
assign OE_DATA_85_const_net_13             = 4'h0;
assign OE_DATA_86_const_net_13             = 4'h0;
assign OE_DATA_87_const_net_13             = 4'h0;
assign OE_DATA_88_const_net_13             = 4'h0;
assign OE_DATA_89_const_net_13             = 4'h0;
assign OE_DATA_90_const_net_13             = 4'h0;
assign OE_DATA_91_const_net_13             = 4'h0;
assign OE_DATA_92_const_net_13             = 4'h0;
assign OE_DATA_93_const_net_13             = 4'h0;
assign OE_DATA_94_const_net_13             = 4'h0;
assign OE_DATA_95_const_net_13             = 4'h0;
assign OE_DATA_96_const_net_13             = 4'h0;
assign OE_DATA_97_const_net_13             = 4'h0;
assign OE_DATA_98_const_net_13             = 4'h0;
assign OE_DATA_99_const_net_13             = 4'h0;
assign OE_DATA_100_const_net_13            = 4'h0;
assign OE_DATA_101_const_net_13            = 4'h0;
assign OE_DATA_102_const_net_13            = 4'h0;
assign OE_DATA_103_const_net_13            = 4'h0;
assign OE_DATA_104_const_net_13            = 4'h0;
assign OE_DATA_105_const_net_13            = 4'h0;
assign OE_DATA_106_const_net_13            = 4'h0;
assign OE_DATA_107_const_net_13            = 4'h0;
assign OE_DATA_108_const_net_13            = 4'h0;
assign OE_DATA_109_const_net_13            = 4'h0;
assign OE_DATA_110_const_net_13            = 4'h0;
assign OE_DATA_111_const_net_13            = 4'h0;
assign OE_DATA_112_const_net_13            = 4'h0;
assign OE_DATA_113_const_net_13            = 4'h0;
assign OE_DATA_114_const_net_13            = 4'h0;
assign OE_DATA_115_const_net_13            = 4'h0;
assign OE_DATA_116_const_net_13            = 4'h0;
assign OE_DATA_117_const_net_13            = 4'h0;
assign OE_DATA_118_const_net_13            = 4'h0;
assign OE_DATA_119_const_net_13            = 4'h0;
assign OE_DATA_120_const_net_13            = 4'h0;
assign OE_DATA_121_const_net_13            = 4'h0;
assign OE_DATA_122_const_net_13            = 4'h0;
assign OE_DATA_123_const_net_13            = 4'h0;
assign OE_DATA_124_const_net_13            = 4'h0;
assign OE_DATA_125_const_net_13            = 4'h0;
assign OE_DATA_126_const_net_13            = 4'h0;
assign OE_DATA_127_const_net_13            = 4'h0;
assign RX_DQS_90_const_net_14              = 2'h0;
assign FIFO_WR_PTR_const_net_14            = 3'h0;
assign FIFO_RD_PTR_const_net_14            = 3'h0;
assign EYE_MONITOR_LANE_WIDTH_const_net_14 = 3'h0;
assign TX_DATA_1_const_net_11              = 4'h0;
assign TX_DATA_2_const_net_13              = 4'h0;
assign TX_DATA_3_const_net_13              = 4'h0;
assign TX_DATA_4_const_net_13              = 4'h0;
assign TX_DATA_5_const_net_13              = 4'h0;
assign TX_DATA_6_const_net_13              = 4'h0;
assign TX_DATA_7_const_net_13              = 4'h0;
assign TX_DATA_8_const_net_13              = 4'h0;
assign TX_DATA_9_const_net_13              = 4'h0;
assign TX_DATA_10_const_net_13             = 4'h0;
assign TX_DATA_11_const_net_13             = 4'h0;
assign TX_DATA_12_const_net_14             = 4'h0;
assign TX_DATA_13_const_net_14             = 4'h0;
assign TX_DATA_14_const_net_14             = 4'h0;
assign TX_DATA_15_const_net_14             = 4'h0;
assign TX_DATA_16_const_net_14             = 4'h0;
assign TX_DATA_17_const_net_14             = 4'h0;
assign TX_DATA_18_const_net_14             = 4'h0;
assign TX_DATA_19_const_net_14             = 4'h0;
assign TX_DATA_20_const_net_14             = 4'h0;
assign TX_DATA_21_const_net_14             = 4'h0;
assign TX_DATA_22_const_net_14             = 4'h0;
assign TX_DATA_23_const_net_14             = 4'h0;
assign TX_DATA_24_const_net_14             = 4'h0;
assign TX_DATA_25_const_net_14             = 4'h0;
assign TX_DATA_26_const_net_14             = 4'h0;
assign TX_DATA_27_const_net_14             = 4'h0;
assign TX_DATA_28_const_net_14             = 4'h0;
assign TX_DATA_29_const_net_14             = 4'h0;
assign TX_DATA_30_const_net_14             = 4'h0;
assign TX_DATA_31_const_net_14             = 4'h0;
assign TX_DATA_32_const_net_14             = 4'h0;
assign TX_DATA_33_const_net_14             = 4'h0;
assign TX_DATA_34_const_net_14             = 4'h0;
assign TX_DATA_35_const_net_14             = 4'h0;
assign TX_DATA_36_const_net_14             = 4'h0;
assign TX_DATA_37_const_net_14             = 4'h0;
assign TX_DATA_38_const_net_14             = 4'h0;
assign TX_DATA_39_const_net_14             = 4'h0;
assign TX_DATA_40_const_net_14             = 4'h0;
assign TX_DATA_41_const_net_14             = 4'h0;
assign TX_DATA_42_const_net_14             = 4'h0;
assign TX_DATA_43_const_net_14             = 4'h0;
assign TX_DATA_44_const_net_14             = 4'h0;
assign TX_DATA_45_const_net_14             = 4'h0;
assign TX_DATA_46_const_net_14             = 4'h0;
assign TX_DATA_47_const_net_14             = 4'h0;
assign TX_DATA_48_const_net_14             = 4'h0;
assign TX_DATA_49_const_net_14             = 4'h0;
assign TX_DATA_50_const_net_14             = 4'h0;
assign TX_DATA_51_const_net_14             = 4'h0;
assign TX_DATA_52_const_net_14             = 4'h0;
assign TX_DATA_53_const_net_14             = 4'h0;
assign TX_DATA_54_const_net_14             = 4'h0;
assign TX_DATA_55_const_net_14             = 4'h0;
assign TX_DATA_56_const_net_14             = 4'h0;
assign TX_DATA_57_const_net_14             = 4'h0;
assign TX_DATA_58_const_net_14             = 4'h0;
assign TX_DATA_59_const_net_14             = 4'h0;
assign TX_DATA_60_const_net_14             = 4'h0;
assign TX_DATA_61_const_net_14             = 4'h0;
assign TX_DATA_62_const_net_14             = 4'h0;
assign TX_DATA_63_const_net_14             = 4'h0;
assign TX_DATA_64_const_net_14             = 4'h0;
assign TX_DATA_65_const_net_14             = 4'h0;
assign TX_DATA_66_const_net_14             = 4'h0;
assign TX_DATA_67_const_net_14             = 4'h0;
assign TX_DATA_68_const_net_14             = 4'h0;
assign TX_DATA_69_const_net_14             = 4'h0;
assign TX_DATA_70_const_net_14             = 4'h0;
assign TX_DATA_71_const_net_14             = 4'h0;
assign TX_DATA_72_const_net_14             = 4'h0;
assign TX_DATA_73_const_net_14             = 4'h0;
assign TX_DATA_74_const_net_14             = 4'h0;
assign TX_DATA_75_const_net_14             = 4'h0;
assign TX_DATA_76_const_net_14             = 4'h0;
assign TX_DATA_77_const_net_14             = 4'h0;
assign TX_DATA_78_const_net_14             = 4'h0;
assign TX_DATA_79_const_net_14             = 4'h0;
assign TX_DATA_80_const_net_14             = 4'h0;
assign TX_DATA_81_const_net_14             = 4'h0;
assign TX_DATA_82_const_net_14             = 4'h0;
assign TX_DATA_83_const_net_14             = 4'h0;
assign TX_DATA_84_const_net_14             = 4'h0;
assign TX_DATA_85_const_net_14             = 4'h0;
assign TX_DATA_86_const_net_14             = 4'h0;
assign TX_DATA_87_const_net_14             = 4'h0;
assign TX_DATA_88_const_net_14             = 4'h0;
assign TX_DATA_89_const_net_14             = 4'h0;
assign TX_DATA_90_const_net_14             = 4'h0;
assign TX_DATA_91_const_net_14             = 4'h0;
assign TX_DATA_92_const_net_14             = 4'h0;
assign TX_DATA_93_const_net_14             = 4'h0;
assign TX_DATA_94_const_net_14             = 4'h0;
assign TX_DATA_95_const_net_14             = 4'h0;
assign TX_DATA_96_const_net_14             = 4'h0;
assign TX_DATA_97_const_net_14             = 4'h0;
assign TX_DATA_98_const_net_14             = 4'h0;
assign TX_DATA_99_const_net_14             = 4'h0;
assign TX_DATA_100_const_net_14            = 4'h0;
assign TX_DATA_101_const_net_14            = 4'h0;
assign TX_DATA_102_const_net_14            = 4'h0;
assign TX_DATA_103_const_net_14            = 4'h0;
assign TX_DATA_104_const_net_14            = 4'h0;
assign TX_DATA_105_const_net_14            = 4'h0;
assign TX_DATA_106_const_net_14            = 4'h0;
assign TX_DATA_107_const_net_14            = 4'h0;
assign TX_DATA_108_const_net_14            = 4'h0;
assign TX_DATA_109_const_net_14            = 4'h0;
assign TX_DATA_110_const_net_14            = 4'h0;
assign TX_DATA_111_const_net_14            = 4'h0;
assign TX_DATA_112_const_net_14            = 4'h0;
assign TX_DATA_113_const_net_14            = 4'h0;
assign TX_DATA_114_const_net_14            = 4'h0;
assign TX_DATA_115_const_net_14            = 4'h0;
assign TX_DATA_116_const_net_14            = 4'h0;
assign TX_DATA_117_const_net_14            = 4'h0;
assign TX_DATA_118_const_net_14            = 4'h0;
assign TX_DATA_119_const_net_14            = 4'h0;
assign TX_DATA_120_const_net_14            = 4'h0;
assign TX_DATA_121_const_net_14            = 4'h0;
assign TX_DATA_122_const_net_14            = 4'h0;
assign TX_DATA_123_const_net_14            = 4'h0;
assign TX_DATA_124_const_net_14            = 4'h0;
assign TX_DATA_125_const_net_14            = 4'h0;
assign TX_DATA_126_const_net_14            = 4'h0;
assign TX_DATA_127_const_net_14            = 4'h0;
assign OE_DATA_1_const_net_14              = 4'h0;
assign OE_DATA_2_const_net_14              = 4'h0;
assign OE_DATA_3_const_net_14              = 4'h0;
assign OE_DATA_4_const_net_14              = 4'h0;
assign OE_DATA_5_const_net_14              = 4'h0;
assign OE_DATA_6_const_net_14              = 4'h0;
assign OE_DATA_7_const_net_14              = 4'h0;
assign OE_DATA_8_const_net_14              = 4'h0;
assign OE_DATA_9_const_net_14              = 4'h0;
assign OE_DATA_10_const_net_14             = 4'h0;
assign OE_DATA_11_const_net_14             = 4'h0;
assign OE_DATA_12_const_net_14             = 4'h0;
assign OE_DATA_13_const_net_14             = 4'h0;
assign OE_DATA_14_const_net_14             = 4'h0;
assign OE_DATA_15_const_net_14             = 4'h0;
assign OE_DATA_16_const_net_14             = 4'h0;
assign OE_DATA_17_const_net_14             = 4'h0;
assign OE_DATA_18_const_net_14             = 4'h0;
assign OE_DATA_19_const_net_14             = 4'h0;
assign OE_DATA_20_const_net_14             = 4'h0;
assign OE_DATA_21_const_net_14             = 4'h0;
assign OE_DATA_22_const_net_14             = 4'h0;
assign OE_DATA_23_const_net_14             = 4'h0;
assign OE_DATA_24_const_net_14             = 4'h0;
assign OE_DATA_25_const_net_14             = 4'h0;
assign OE_DATA_26_const_net_14             = 4'h0;
assign OE_DATA_27_const_net_14             = 4'h0;
assign OE_DATA_28_const_net_14             = 4'h0;
assign OE_DATA_29_const_net_14             = 4'h0;
assign OE_DATA_30_const_net_14             = 4'h0;
assign OE_DATA_31_const_net_14             = 4'h0;
assign OE_DATA_32_const_net_14             = 4'h0;
assign OE_DATA_33_const_net_14             = 4'h0;
assign OE_DATA_34_const_net_14             = 4'h0;
assign OE_DATA_35_const_net_14             = 4'h0;
assign OE_DATA_36_const_net_14             = 4'h0;
assign OE_DATA_37_const_net_14             = 4'h0;
assign OE_DATA_38_const_net_14             = 4'h0;
assign OE_DATA_39_const_net_14             = 4'h0;
assign OE_DATA_40_const_net_14             = 4'h0;
assign OE_DATA_41_const_net_14             = 4'h0;
assign OE_DATA_42_const_net_14             = 4'h0;
assign OE_DATA_43_const_net_14             = 4'h0;
assign OE_DATA_44_const_net_14             = 4'h0;
assign OE_DATA_45_const_net_14             = 4'h0;
assign OE_DATA_46_const_net_14             = 4'h0;
assign OE_DATA_47_const_net_14             = 4'h0;
assign OE_DATA_48_const_net_14             = 4'h0;
assign OE_DATA_49_const_net_14             = 4'h0;
assign OE_DATA_50_const_net_14             = 4'h0;
assign OE_DATA_51_const_net_14             = 4'h0;
assign OE_DATA_52_const_net_14             = 4'h0;
assign OE_DATA_53_const_net_14             = 4'h0;
assign OE_DATA_54_const_net_14             = 4'h0;
assign OE_DATA_55_const_net_14             = 4'h0;
assign OE_DATA_56_const_net_14             = 4'h0;
assign OE_DATA_57_const_net_14             = 4'h0;
assign OE_DATA_58_const_net_14             = 4'h0;
assign OE_DATA_59_const_net_14             = 4'h0;
assign OE_DATA_60_const_net_14             = 4'h0;
assign OE_DATA_61_const_net_14             = 4'h0;
assign OE_DATA_62_const_net_14             = 4'h0;
assign OE_DATA_63_const_net_14             = 4'h0;
assign OE_DATA_64_const_net_14             = 4'h0;
assign OE_DATA_65_const_net_14             = 4'h0;
assign OE_DATA_66_const_net_14             = 4'h0;
assign OE_DATA_67_const_net_14             = 4'h0;
assign OE_DATA_68_const_net_14             = 4'h0;
assign OE_DATA_69_const_net_14             = 4'h0;
assign OE_DATA_70_const_net_14             = 4'h0;
assign OE_DATA_71_const_net_14             = 4'h0;
assign OE_DATA_72_const_net_14             = 4'h0;
assign OE_DATA_73_const_net_14             = 4'h0;
assign OE_DATA_74_const_net_14             = 4'h0;
assign OE_DATA_75_const_net_14             = 4'h0;
assign OE_DATA_76_const_net_14             = 4'h0;
assign OE_DATA_77_const_net_14             = 4'h0;
assign OE_DATA_78_const_net_14             = 4'h0;
assign OE_DATA_79_const_net_14             = 4'h0;
assign OE_DATA_80_const_net_14             = 4'h0;
assign OE_DATA_81_const_net_14             = 4'h0;
assign OE_DATA_82_const_net_14             = 4'h0;
assign OE_DATA_83_const_net_14             = 4'h0;
assign OE_DATA_84_const_net_14             = 4'h0;
assign OE_DATA_85_const_net_14             = 4'h0;
assign OE_DATA_86_const_net_14             = 4'h0;
assign OE_DATA_87_const_net_14             = 4'h0;
assign OE_DATA_88_const_net_14             = 4'h0;
assign OE_DATA_89_const_net_14             = 4'h0;
assign OE_DATA_90_const_net_14             = 4'h0;
assign OE_DATA_91_const_net_14             = 4'h0;
assign OE_DATA_92_const_net_14             = 4'h0;
assign OE_DATA_93_const_net_14             = 4'h0;
assign OE_DATA_94_const_net_14             = 4'h0;
assign OE_DATA_95_const_net_14             = 4'h0;
assign OE_DATA_96_const_net_14             = 4'h0;
assign OE_DATA_97_const_net_14             = 4'h0;
assign OE_DATA_98_const_net_14             = 4'h0;
assign OE_DATA_99_const_net_14             = 4'h0;
assign OE_DATA_100_const_net_14            = 4'h0;
assign OE_DATA_101_const_net_14            = 4'h0;
assign OE_DATA_102_const_net_14            = 4'h0;
assign OE_DATA_103_const_net_14            = 4'h0;
assign OE_DATA_104_const_net_14            = 4'h0;
assign OE_DATA_105_const_net_14            = 4'h0;
assign OE_DATA_106_const_net_14            = 4'h0;
assign OE_DATA_107_const_net_14            = 4'h0;
assign OE_DATA_108_const_net_14            = 4'h0;
assign OE_DATA_109_const_net_14            = 4'h0;
assign OE_DATA_110_const_net_14            = 4'h0;
assign OE_DATA_111_const_net_14            = 4'h0;
assign OE_DATA_112_const_net_14            = 4'h0;
assign OE_DATA_113_const_net_14            = 4'h0;
assign OE_DATA_114_const_net_14            = 4'h0;
assign OE_DATA_115_const_net_14            = 4'h0;
assign OE_DATA_116_const_net_14            = 4'h0;
assign OE_DATA_117_const_net_14            = 4'h0;
assign OE_DATA_118_const_net_14            = 4'h0;
assign OE_DATA_119_const_net_14            = 4'h0;
assign OE_DATA_120_const_net_14            = 4'h0;
assign OE_DATA_121_const_net_14            = 4'h0;
assign OE_DATA_122_const_net_14            = 4'h0;
assign OE_DATA_123_const_net_14            = 4'h0;
assign OE_DATA_124_const_net_14            = 4'h0;
assign OE_DATA_125_const_net_14            = 4'h0;
assign OE_DATA_126_const_net_14            = 4'h0;
assign OE_DATA_127_const_net_14            = 4'h0;
assign CDR_CLK_B_SEL_const_net_0           = 11'h000;
assign FIFO_WR_PTR_const_net_15            = 3'h0;
assign FIFO_RD_PTR_const_net_15            = 3'h0;
assign EYE_MONITOR_LANE_WIDTH_const_net_15 = 3'h0;
assign TX_DATA_1_const_net_12              = 8'h00;
assign TX_DATA_2_const_net_14              = 8'h00;
assign TX_DATA_3_const_net_14              = 8'h00;
assign TX_DATA_4_const_net_14              = 8'h00;
assign TX_DATA_5_const_net_14              = 8'h00;
assign TX_DATA_6_const_net_14              = 8'h00;
assign TX_DATA_7_const_net_14              = 8'h00;
assign TX_DATA_8_const_net_14              = 8'h00;
assign TX_DATA_9_const_net_14              = 8'h00;
assign TX_DATA_10_const_net_14             = 8'h00;
assign TX_DATA_11_const_net_14             = 8'h00;
assign TX_DATA_12_const_net_15             = 8'h00;
assign TX_DATA_13_const_net_15             = 8'h00;
assign TX_DATA_14_const_net_15             = 8'h00;
assign TX_DATA_15_const_net_15             = 8'h00;
assign TX_DATA_16_const_net_15             = 8'h00;
assign TX_DATA_17_const_net_15             = 8'h00;
assign TX_DATA_18_const_net_15             = 8'h00;
assign TX_DATA_19_const_net_15             = 8'h00;
assign TX_DATA_20_const_net_15             = 8'h00;
assign TX_DATA_21_const_net_15             = 8'h00;
assign TX_DATA_22_const_net_15             = 8'h00;
assign TX_DATA_23_const_net_15             = 8'h00;
assign TX_DATA_24_const_net_15             = 8'h00;
assign TX_DATA_25_const_net_15             = 8'h00;
assign TX_DATA_26_const_net_15             = 8'h00;
assign TX_DATA_27_const_net_15             = 8'h00;
assign TX_DATA_28_const_net_15             = 8'h00;
assign TX_DATA_29_const_net_15             = 8'h00;
assign TX_DATA_30_const_net_15             = 8'h00;
assign TX_DATA_31_const_net_15             = 8'h00;
assign TX_DATA_32_const_net_15             = 8'h00;
assign TX_DATA_33_const_net_15             = 8'h00;
assign TX_DATA_34_const_net_15             = 8'h00;
assign TX_DATA_35_const_net_15             = 8'h00;
assign TX_DATA_36_const_net_15             = 8'h00;
assign TX_DATA_37_const_net_15             = 8'h00;
assign TX_DATA_38_const_net_15             = 8'h00;
assign TX_DATA_39_const_net_15             = 8'h00;
assign TX_DATA_40_const_net_15             = 8'h00;
assign TX_DATA_41_const_net_15             = 8'h00;
assign TX_DATA_42_const_net_15             = 8'h00;
assign TX_DATA_43_const_net_15             = 8'h00;
assign TX_DATA_44_const_net_15             = 8'h00;
assign TX_DATA_45_const_net_15             = 8'h00;
assign TX_DATA_46_const_net_15             = 8'h00;
assign TX_DATA_47_const_net_15             = 8'h00;
assign TX_DATA_48_const_net_15             = 8'h00;
assign TX_DATA_49_const_net_15             = 8'h00;
assign TX_DATA_50_const_net_15             = 8'h00;
assign TX_DATA_51_const_net_15             = 8'h00;
assign TX_DATA_52_const_net_15             = 8'h00;
assign TX_DATA_53_const_net_15             = 8'h00;
assign TX_DATA_54_const_net_15             = 8'h00;
assign TX_DATA_55_const_net_15             = 8'h00;
assign TX_DATA_56_const_net_15             = 8'h00;
assign TX_DATA_57_const_net_15             = 8'h00;
assign TX_DATA_58_const_net_15             = 8'h00;
assign TX_DATA_59_const_net_15             = 8'h00;
assign TX_DATA_60_const_net_15             = 8'h00;
assign TX_DATA_61_const_net_15             = 8'h00;
assign TX_DATA_62_const_net_15             = 8'h00;
assign TX_DATA_63_const_net_15             = 8'h00;
assign TX_DATA_64_const_net_15             = 8'h00;
assign TX_DATA_65_const_net_15             = 8'h00;
assign TX_DATA_66_const_net_15             = 8'h00;
assign TX_DATA_67_const_net_15             = 8'h00;
assign TX_DATA_68_const_net_15             = 8'h00;
assign TX_DATA_69_const_net_15             = 8'h00;
assign TX_DATA_70_const_net_15             = 8'h00;
assign TX_DATA_71_const_net_15             = 8'h00;
assign TX_DATA_72_const_net_15             = 8'h00;
assign TX_DATA_73_const_net_15             = 8'h00;
assign TX_DATA_74_const_net_15             = 8'h00;
assign TX_DATA_75_const_net_15             = 8'h00;
assign TX_DATA_76_const_net_15             = 8'h00;
assign TX_DATA_77_const_net_15             = 8'h00;
assign TX_DATA_78_const_net_15             = 8'h00;
assign TX_DATA_79_const_net_15             = 8'h00;
assign TX_DATA_80_const_net_15             = 8'h00;
assign TX_DATA_81_const_net_15             = 8'h00;
assign TX_DATA_82_const_net_15             = 8'h00;
assign TX_DATA_83_const_net_15             = 8'h00;
assign TX_DATA_84_const_net_15             = 8'h00;
assign TX_DATA_85_const_net_15             = 8'h00;
assign TX_DATA_86_const_net_15             = 8'h00;
assign TX_DATA_87_const_net_15             = 8'h00;
assign TX_DATA_88_const_net_15             = 8'h00;
assign TX_DATA_89_const_net_15             = 8'h00;
assign TX_DATA_90_const_net_15             = 8'h00;
assign TX_DATA_91_const_net_15             = 8'h00;
assign TX_DATA_92_const_net_15             = 8'h00;
assign TX_DATA_93_const_net_15             = 8'h00;
assign TX_DATA_94_const_net_15             = 8'h00;
assign TX_DATA_95_const_net_15             = 8'h00;
assign TX_DATA_96_const_net_15             = 8'h00;
assign TX_DATA_97_const_net_15             = 8'h00;
assign TX_DATA_98_const_net_15             = 8'h00;
assign TX_DATA_99_const_net_15             = 8'h00;
assign TX_DATA_100_const_net_15            = 8'h00;
assign TX_DATA_101_const_net_15            = 8'h00;
assign TX_DATA_102_const_net_15            = 8'h00;
assign TX_DATA_103_const_net_15            = 8'h00;
assign TX_DATA_104_const_net_15            = 8'h00;
assign TX_DATA_105_const_net_15            = 8'h00;
assign TX_DATA_106_const_net_15            = 8'h00;
assign TX_DATA_107_const_net_15            = 8'h00;
assign TX_DATA_108_const_net_15            = 8'h00;
assign TX_DATA_109_const_net_15            = 8'h00;
assign TX_DATA_110_const_net_15            = 8'h00;
assign TX_DATA_111_const_net_15            = 8'h00;
assign TX_DATA_112_const_net_15            = 8'h00;
assign TX_DATA_113_const_net_15            = 8'h00;
assign TX_DATA_114_const_net_15            = 8'h00;
assign TX_DATA_115_const_net_15            = 8'h00;
assign TX_DATA_116_const_net_15            = 8'h00;
assign TX_DATA_117_const_net_15            = 8'h00;
assign TX_DATA_118_const_net_15            = 8'h00;
assign TX_DATA_119_const_net_15            = 8'h00;
assign TX_DATA_120_const_net_15            = 8'h00;
assign TX_DATA_121_const_net_15            = 8'h00;
assign TX_DATA_122_const_net_15            = 8'h00;
assign TX_DATA_123_const_net_15            = 8'h00;
assign TX_DATA_124_const_net_15            = 8'h00;
assign TX_DATA_125_const_net_15            = 8'h00;
assign TX_DATA_126_const_net_15            = 8'h00;
assign TX_DATA_127_const_net_15            = 8'h00;
assign OE_DATA_1_const_net_15              = 4'h0;
assign OE_DATA_2_const_net_15              = 4'h0;
assign OE_DATA_3_const_net_15              = 4'h0;
assign OE_DATA_4_const_net_15              = 4'h0;
assign OE_DATA_5_const_net_15              = 4'h0;
assign OE_DATA_6_const_net_15              = 4'h0;
assign OE_DATA_7_const_net_15              = 4'h0;
assign OE_DATA_8_const_net_15              = 4'h0;
assign OE_DATA_9_const_net_15              = 4'h0;
assign OE_DATA_10_const_net_15             = 4'h0;
assign OE_DATA_11_const_net_15             = 4'h0;
assign OE_DATA_12_const_net_15             = 4'h0;
assign OE_DATA_13_const_net_15             = 4'h0;
assign OE_DATA_14_const_net_15             = 4'h0;
assign OE_DATA_15_const_net_15             = 4'h0;
assign OE_DATA_16_const_net_15             = 4'h0;
assign OE_DATA_17_const_net_15             = 4'h0;
assign OE_DATA_18_const_net_15             = 4'h0;
assign OE_DATA_19_const_net_15             = 4'h0;
assign OE_DATA_20_const_net_15             = 4'h0;
assign OE_DATA_21_const_net_15             = 4'h0;
assign OE_DATA_22_const_net_15             = 4'h0;
assign OE_DATA_23_const_net_15             = 4'h0;
assign OE_DATA_24_const_net_15             = 4'h0;
assign OE_DATA_25_const_net_15             = 4'h0;
assign OE_DATA_26_const_net_15             = 4'h0;
assign OE_DATA_27_const_net_15             = 4'h0;
assign OE_DATA_28_const_net_15             = 4'h0;
assign OE_DATA_29_const_net_15             = 4'h0;
assign OE_DATA_30_const_net_15             = 4'h0;
assign OE_DATA_31_const_net_15             = 4'h0;
assign OE_DATA_32_const_net_15             = 4'h0;
assign OE_DATA_33_const_net_15             = 4'h0;
assign OE_DATA_34_const_net_15             = 4'h0;
assign OE_DATA_35_const_net_15             = 4'h0;
assign OE_DATA_36_const_net_15             = 4'h0;
assign OE_DATA_37_const_net_15             = 4'h0;
assign OE_DATA_38_const_net_15             = 4'h0;
assign OE_DATA_39_const_net_15             = 4'h0;
assign OE_DATA_40_const_net_15             = 4'h0;
assign OE_DATA_41_const_net_15             = 4'h0;
assign OE_DATA_42_const_net_15             = 4'h0;
assign OE_DATA_43_const_net_15             = 4'h0;
assign OE_DATA_44_const_net_15             = 4'h0;
assign OE_DATA_45_const_net_15             = 4'h0;
assign OE_DATA_46_const_net_15             = 4'h0;
assign OE_DATA_47_const_net_15             = 4'h0;
assign OE_DATA_48_const_net_15             = 4'h0;
assign OE_DATA_49_const_net_15             = 4'h0;
assign OE_DATA_50_const_net_15             = 4'h0;
assign OE_DATA_51_const_net_15             = 4'h0;
assign OE_DATA_52_const_net_15             = 4'h0;
assign OE_DATA_53_const_net_15             = 4'h0;
assign OE_DATA_54_const_net_15             = 4'h0;
assign OE_DATA_55_const_net_15             = 4'h0;
assign OE_DATA_56_const_net_15             = 4'h0;
assign OE_DATA_57_const_net_15             = 4'h0;
assign OE_DATA_58_const_net_15             = 4'h0;
assign OE_DATA_59_const_net_15             = 4'h0;
assign OE_DATA_60_const_net_15             = 4'h0;
assign OE_DATA_61_const_net_15             = 4'h0;
assign OE_DATA_62_const_net_15             = 4'h0;
assign OE_DATA_63_const_net_15             = 4'h0;
assign OE_DATA_64_const_net_15             = 4'h0;
assign OE_DATA_65_const_net_15             = 4'h0;
assign OE_DATA_66_const_net_15             = 4'h0;
assign OE_DATA_67_const_net_15             = 4'h0;
assign OE_DATA_68_const_net_15             = 4'h0;
assign OE_DATA_69_const_net_15             = 4'h0;
assign OE_DATA_70_const_net_15             = 4'h0;
assign OE_DATA_71_const_net_15             = 4'h0;
assign OE_DATA_72_const_net_15             = 4'h0;
assign OE_DATA_73_const_net_15             = 4'h0;
assign OE_DATA_74_const_net_15             = 4'h0;
assign OE_DATA_75_const_net_15             = 4'h0;
assign OE_DATA_76_const_net_15             = 4'h0;
assign OE_DATA_77_const_net_15             = 4'h0;
assign OE_DATA_78_const_net_15             = 4'h0;
assign OE_DATA_79_const_net_15             = 4'h0;
assign OE_DATA_80_const_net_15             = 4'h0;
assign OE_DATA_81_const_net_15             = 4'h0;
assign OE_DATA_82_const_net_15             = 4'h0;
assign OE_DATA_83_const_net_15             = 4'h0;
assign OE_DATA_84_const_net_15             = 4'h0;
assign OE_DATA_85_const_net_15             = 4'h0;
assign OE_DATA_86_const_net_15             = 4'h0;
assign OE_DATA_87_const_net_15             = 4'h0;
assign OE_DATA_88_const_net_15             = 4'h0;
assign OE_DATA_89_const_net_15             = 4'h0;
assign OE_DATA_90_const_net_15             = 4'h0;
assign OE_DATA_91_const_net_15             = 4'h0;
assign OE_DATA_92_const_net_15             = 4'h0;
assign OE_DATA_93_const_net_15             = 4'h0;
assign OE_DATA_94_const_net_15             = 4'h0;
assign OE_DATA_95_const_net_15             = 4'h0;
assign OE_DATA_96_const_net_15             = 4'h0;
assign OE_DATA_97_const_net_15             = 4'h0;
assign OE_DATA_98_const_net_15             = 4'h0;
assign OE_DATA_99_const_net_15             = 4'h0;
assign OE_DATA_100_const_net_15            = 4'h0;
assign OE_DATA_101_const_net_15            = 4'h0;
assign OE_DATA_102_const_net_15            = 4'h0;
assign OE_DATA_103_const_net_15            = 4'h0;
assign OE_DATA_104_const_net_15            = 4'h0;
assign OE_DATA_105_const_net_15            = 4'h0;
assign OE_DATA_106_const_net_15            = 4'h0;
assign OE_DATA_107_const_net_15            = 4'h0;
assign OE_DATA_108_const_net_15            = 4'h0;
assign OE_DATA_109_const_net_15            = 4'h0;
assign OE_DATA_110_const_net_15            = 4'h0;
assign OE_DATA_111_const_net_15            = 4'h0;
assign OE_DATA_112_const_net_15            = 4'h0;
assign OE_DATA_113_const_net_15            = 4'h0;
assign OE_DATA_114_const_net_15            = 4'h0;
assign OE_DATA_115_const_net_15            = 4'h0;
assign OE_DATA_116_const_net_15            = 4'h0;
assign OE_DATA_117_const_net_15            = 4'h0;
assign OE_DATA_118_const_net_15            = 4'h0;
assign OE_DATA_119_const_net_15            = 4'h0;
assign OE_DATA_120_const_net_15            = 4'h0;
assign OE_DATA_121_const_net_15            = 4'h0;
assign OE_DATA_122_const_net_15            = 4'h0;
assign OE_DATA_123_const_net_15            = 4'h0;
assign OE_DATA_124_const_net_15            = 4'h0;
assign OE_DATA_125_const_net_15            = 4'h0;
assign OE_DATA_126_const_net_15            = 4'h0;
assign OE_DATA_127_const_net_15            = 4'h0;
assign TX_DATA_8_const_net_15              = 8'h00;
assign TX_DATA_9_const_net_15              = 8'h00;
assign TX_DATA_10_const_net_15             = 8'h00;
assign TX_DATA_11_const_net_15             = 8'h00;
assign TX_DATA_12_const_net_16             = 8'h00;
assign TX_DATA_13_const_net_16             = 8'h00;
assign TX_DATA_14_const_net_16             = 8'h00;
assign TX_DATA_15_const_net_16             = 8'h00;
assign TX_DATA_16_const_net_16             = 8'h00;
assign TX_DATA_17_const_net_16             = 8'h00;
assign TX_DATA_18_const_net_16             = 8'h00;
assign TX_DATA_19_const_net_16             = 8'h00;
assign TX_DATA_20_const_net_16             = 8'h00;
assign TX_DATA_21_const_net_16             = 8'h00;
assign TX_DATA_22_const_net_16             = 8'h00;
assign TX_DATA_23_const_net_16             = 8'h00;
assign TX_DATA_24_const_net_16             = 8'h00;
assign TX_DATA_25_const_net_16             = 8'h00;
assign TX_DATA_26_const_net_16             = 8'h00;
assign TX_DATA_27_const_net_16             = 8'h00;
assign TX_DATA_28_const_net_16             = 8'h00;
assign TX_DATA_29_const_net_16             = 8'h00;
assign TX_DATA_30_const_net_16             = 8'h00;
assign TX_DATA_31_const_net_16             = 8'h00;
assign TX_DATA_32_const_net_16             = 8'h00;
assign TX_DATA_33_const_net_16             = 8'h00;
assign TX_DATA_34_const_net_16             = 8'h00;
assign TX_DATA_35_const_net_16             = 8'h00;
assign TX_DATA_36_const_net_16             = 8'h00;
assign TX_DATA_37_const_net_16             = 8'h00;
assign TX_DATA_38_const_net_16             = 8'h00;
assign TX_DATA_39_const_net_16             = 8'h00;
assign TX_DATA_40_const_net_16             = 8'h00;
assign TX_DATA_41_const_net_16             = 8'h00;
assign TX_DATA_42_const_net_16             = 8'h00;
assign TX_DATA_43_const_net_16             = 8'h00;
assign TX_DATA_44_const_net_16             = 8'h00;
assign TX_DATA_45_const_net_16             = 8'h00;
assign TX_DATA_46_const_net_16             = 8'h00;
assign TX_DATA_47_const_net_16             = 8'h00;
assign TX_DATA_48_const_net_16             = 8'h00;
assign TX_DATA_49_const_net_16             = 8'h00;
assign TX_DATA_50_const_net_16             = 8'h00;
assign TX_DATA_51_const_net_16             = 8'h00;
assign TX_DATA_52_const_net_16             = 8'h00;
assign TX_DATA_53_const_net_16             = 8'h00;
assign TX_DATA_54_const_net_16             = 8'h00;
assign TX_DATA_55_const_net_16             = 8'h00;
assign TX_DATA_56_const_net_16             = 8'h00;
assign TX_DATA_57_const_net_16             = 8'h00;
assign TX_DATA_58_const_net_16             = 8'h00;
assign TX_DATA_59_const_net_16             = 8'h00;
assign TX_DATA_60_const_net_16             = 8'h00;
assign TX_DATA_61_const_net_16             = 8'h00;
assign TX_DATA_62_const_net_16             = 8'h00;
assign TX_DATA_63_const_net_16             = 8'h00;
assign TX_DATA_64_const_net_16             = 8'h00;
assign TX_DATA_65_const_net_16             = 8'h00;
assign TX_DATA_66_const_net_16             = 8'h00;
assign TX_DATA_67_const_net_16             = 8'h00;
assign TX_DATA_68_const_net_16             = 8'h00;
assign TX_DATA_69_const_net_16             = 8'h00;
assign TX_DATA_70_const_net_16             = 8'h00;
assign TX_DATA_71_const_net_16             = 8'h00;
assign TX_DATA_72_const_net_16             = 8'h00;
assign TX_DATA_73_const_net_16             = 8'h00;
assign TX_DATA_74_const_net_16             = 8'h00;
assign TX_DATA_75_const_net_16             = 8'h00;
assign TX_DATA_76_const_net_16             = 8'h00;
assign TX_DATA_77_const_net_16             = 8'h00;
assign TX_DATA_78_const_net_16             = 8'h00;
assign TX_DATA_79_const_net_16             = 8'h00;
assign TX_DATA_80_const_net_16             = 8'h00;
assign TX_DATA_81_const_net_16             = 8'h00;
assign TX_DATA_82_const_net_16             = 8'h00;
assign TX_DATA_83_const_net_16             = 8'h00;
assign TX_DATA_84_const_net_16             = 8'h00;
assign TX_DATA_85_const_net_16             = 8'h00;
assign TX_DATA_86_const_net_16             = 8'h00;
assign TX_DATA_87_const_net_16             = 8'h00;
assign TX_DATA_88_const_net_16             = 8'h00;
assign TX_DATA_89_const_net_16             = 8'h00;
assign TX_DATA_90_const_net_16             = 8'h00;
assign TX_DATA_91_const_net_16             = 8'h00;
assign TX_DATA_92_const_net_16             = 8'h00;
assign TX_DATA_93_const_net_16             = 8'h00;
assign TX_DATA_94_const_net_16             = 8'h00;
assign TX_DATA_95_const_net_16             = 8'h00;
assign TX_DATA_96_const_net_16             = 8'h00;
assign TX_DATA_97_const_net_16             = 8'h00;
assign TX_DATA_98_const_net_16             = 8'h00;
assign TX_DATA_99_const_net_16             = 8'h00;
assign TX_DATA_100_const_net_16            = 8'h00;
assign TX_DATA_101_const_net_16            = 8'h00;
assign TX_DATA_102_const_net_16            = 8'h00;
assign TX_DATA_103_const_net_16            = 8'h00;
assign TX_DATA_104_const_net_16            = 8'h00;
assign TX_DATA_105_const_net_16            = 8'h00;
assign TX_DATA_106_const_net_16            = 8'h00;
assign TX_DATA_107_const_net_16            = 8'h00;
assign TX_DATA_108_const_net_16            = 8'h00;
assign TX_DATA_109_const_net_16            = 8'h00;
assign TX_DATA_110_const_net_16            = 8'h00;
assign TX_DATA_111_const_net_16            = 8'h00;
assign TX_DATA_112_const_net_16            = 8'h00;
assign TX_DATA_113_const_net_16            = 8'h00;
assign TX_DATA_114_const_net_16            = 8'h00;
assign TX_DATA_115_const_net_16            = 8'h00;
assign TX_DATA_116_const_net_16            = 8'h00;
assign TX_DATA_117_const_net_16            = 8'h00;
assign TX_DATA_118_const_net_16            = 8'h00;
assign TX_DATA_119_const_net_16            = 8'h00;
assign TX_DATA_120_const_net_16            = 8'h00;
assign TX_DATA_121_const_net_16            = 8'h00;
assign TX_DATA_122_const_net_16            = 8'h00;
assign TX_DATA_123_const_net_16            = 8'h00;
assign TX_DATA_124_const_net_16            = 8'h00;
assign TX_DATA_125_const_net_16            = 8'h00;
assign TX_DATA_126_const_net_16            = 8'h00;
assign TX_DATA_127_const_net_16            = 8'h00;
assign OE_DATA_8_const_net_16              = 4'h0;
assign OE_DATA_9_const_net_16              = 4'h0;
assign OE_DATA_10_const_net_16             = 4'h0;
assign OE_DATA_11_const_net_16             = 4'h0;
assign OE_DATA_12_const_net_16             = 4'h0;
assign OE_DATA_13_const_net_16             = 4'h0;
assign OE_DATA_14_const_net_16             = 4'h0;
assign OE_DATA_15_const_net_16             = 4'h0;
assign OE_DATA_16_const_net_16             = 4'h0;
assign OE_DATA_17_const_net_16             = 4'h0;
assign OE_DATA_18_const_net_16             = 4'h0;
assign OE_DATA_19_const_net_16             = 4'h0;
assign OE_DATA_20_const_net_16             = 4'h0;
assign OE_DATA_21_const_net_16             = 4'h0;
assign OE_DATA_22_const_net_16             = 4'h0;
assign OE_DATA_23_const_net_16             = 4'h0;
assign OE_DATA_24_const_net_16             = 4'h0;
assign OE_DATA_25_const_net_16             = 4'h0;
assign OE_DATA_26_const_net_16             = 4'h0;
assign OE_DATA_27_const_net_16             = 4'h0;
assign OE_DATA_28_const_net_16             = 4'h0;
assign OE_DATA_29_const_net_16             = 4'h0;
assign OE_DATA_30_const_net_16             = 4'h0;
assign OE_DATA_31_const_net_16             = 4'h0;
assign OE_DATA_32_const_net_16             = 4'h0;
assign OE_DATA_33_const_net_16             = 4'h0;
assign OE_DATA_34_const_net_16             = 4'h0;
assign OE_DATA_35_const_net_16             = 4'h0;
assign OE_DATA_36_const_net_16             = 4'h0;
assign OE_DATA_37_const_net_16             = 4'h0;
assign OE_DATA_38_const_net_16             = 4'h0;
assign OE_DATA_39_const_net_16             = 4'h0;
assign OE_DATA_40_const_net_16             = 4'h0;
assign OE_DATA_41_const_net_16             = 4'h0;
assign OE_DATA_42_const_net_16             = 4'h0;
assign OE_DATA_43_const_net_16             = 4'h0;
assign OE_DATA_44_const_net_16             = 4'h0;
assign OE_DATA_45_const_net_16             = 4'h0;
assign OE_DATA_46_const_net_16             = 4'h0;
assign OE_DATA_47_const_net_16             = 4'h0;
assign OE_DATA_48_const_net_16             = 4'h0;
assign OE_DATA_49_const_net_16             = 4'h0;
assign OE_DATA_50_const_net_16             = 4'h0;
assign OE_DATA_51_const_net_16             = 4'h0;
assign OE_DATA_52_const_net_16             = 4'h0;
assign OE_DATA_53_const_net_16             = 4'h0;
assign OE_DATA_54_const_net_16             = 4'h0;
assign OE_DATA_55_const_net_16             = 4'h0;
assign OE_DATA_56_const_net_16             = 4'h0;
assign OE_DATA_57_const_net_16             = 4'h0;
assign OE_DATA_58_const_net_16             = 4'h0;
assign OE_DATA_59_const_net_16             = 4'h0;
assign OE_DATA_60_const_net_16             = 4'h0;
assign OE_DATA_61_const_net_16             = 4'h0;
assign OE_DATA_62_const_net_16             = 4'h0;
assign OE_DATA_63_const_net_16             = 4'h0;
assign OE_DATA_64_const_net_16             = 4'h0;
assign OE_DATA_65_const_net_16             = 4'h0;
assign OE_DATA_66_const_net_16             = 4'h0;
assign OE_DATA_67_const_net_16             = 4'h0;
assign OE_DATA_68_const_net_16             = 4'h0;
assign OE_DATA_69_const_net_16             = 4'h0;
assign OE_DATA_70_const_net_16             = 4'h0;
assign OE_DATA_71_const_net_16             = 4'h0;
assign OE_DATA_72_const_net_16             = 4'h0;
assign OE_DATA_73_const_net_16             = 4'h0;
assign OE_DATA_74_const_net_16             = 4'h0;
assign OE_DATA_75_const_net_16             = 4'h0;
assign OE_DATA_76_const_net_16             = 4'h0;
assign OE_DATA_77_const_net_16             = 4'h0;
assign OE_DATA_78_const_net_16             = 4'h0;
assign OE_DATA_79_const_net_16             = 4'h0;
assign OE_DATA_80_const_net_16             = 4'h0;
assign OE_DATA_81_const_net_16             = 4'h0;
assign OE_DATA_82_const_net_16             = 4'h0;
assign OE_DATA_83_const_net_16             = 4'h0;
assign OE_DATA_84_const_net_16             = 4'h0;
assign OE_DATA_85_const_net_16             = 4'h0;
assign OE_DATA_86_const_net_16             = 4'h0;
assign OE_DATA_87_const_net_16             = 4'h0;
assign OE_DATA_88_const_net_16             = 4'h0;
assign OE_DATA_89_const_net_16             = 4'h0;
assign OE_DATA_90_const_net_16             = 4'h0;
assign OE_DATA_91_const_net_16             = 4'h0;
assign OE_DATA_92_const_net_16             = 4'h0;
assign OE_DATA_93_const_net_16             = 4'h0;
assign OE_DATA_94_const_net_16             = 4'h0;
assign OE_DATA_95_const_net_16             = 4'h0;
assign OE_DATA_96_const_net_16             = 4'h0;
assign OE_DATA_97_const_net_16             = 4'h0;
assign OE_DATA_98_const_net_16             = 4'h0;
assign OE_DATA_99_const_net_16             = 4'h0;
assign OE_DATA_100_const_net_16            = 4'h0;
assign OE_DATA_101_const_net_16            = 4'h0;
assign OE_DATA_102_const_net_16            = 4'h0;
assign OE_DATA_103_const_net_16            = 4'h0;
assign OE_DATA_104_const_net_16            = 4'h0;
assign OE_DATA_105_const_net_16            = 4'h0;
assign OE_DATA_106_const_net_16            = 4'h0;
assign OE_DATA_107_const_net_16            = 4'h0;
assign OE_DATA_108_const_net_16            = 4'h0;
assign OE_DATA_109_const_net_16            = 4'h0;
assign OE_DATA_110_const_net_16            = 4'h0;
assign OE_DATA_111_const_net_16            = 4'h0;
assign OE_DATA_112_const_net_16            = 4'h0;
assign OE_DATA_113_const_net_16            = 4'h0;
assign OE_DATA_114_const_net_16            = 4'h0;
assign OE_DATA_115_const_net_16            = 4'h0;
assign OE_DATA_116_const_net_16            = 4'h0;
assign OE_DATA_117_const_net_16            = 4'h0;
assign OE_DATA_118_const_net_16            = 4'h0;
assign OE_DATA_119_const_net_16            = 4'h0;
assign OE_DATA_120_const_net_16            = 4'h0;
assign OE_DATA_121_const_net_16            = 4'h0;
assign OE_DATA_122_const_net_16            = 4'h0;
assign OE_DATA_123_const_net_16            = 4'h0;
assign OE_DATA_124_const_net_16            = 4'h0;
assign OE_DATA_125_const_net_16            = 4'h0;
assign OE_DATA_126_const_net_16            = 4'h0;
assign OE_DATA_127_const_net_16            = 4'h0;
assign PAD_I_const_net_3                   = 8'h00;
assign PAD_N_const_net_3                   = 8'h00;
assign PAD_I_N_const_net_3                 = 8'h00;
assign TX_DATA_1_const_net_13              = 8'h00;
assign TX_DATA_2_const_net_15              = 8'h00;
assign TX_DATA_3_const_net_15              = 8'h00;
assign TX_DATA_4_const_net_15              = 8'h00;
assign TX_DATA_5_const_net_15              = 8'h00;
assign TX_DATA_6_const_net_15              = 8'h00;
assign TX_DATA_7_const_net_15              = 8'h00;
assign TX_DATA_8_const_net_16              = 8'h00;
assign TX_DATA_9_const_net_16              = 8'h00;
assign TX_DATA_10_const_net_16             = 8'h00;
assign TX_DATA_11_const_net_16             = 8'h00;
assign TX_DATA_12_const_net_17             = 8'h00;
assign TX_DATA_13_const_net_17             = 8'h00;
assign TX_DATA_14_const_net_17             = 8'h00;
assign TX_DATA_15_const_net_17             = 8'h00;
assign TX_DATA_16_const_net_17             = 8'h00;
assign TX_DATA_17_const_net_17             = 8'h00;
assign TX_DATA_18_const_net_17             = 8'h00;
assign TX_DATA_19_const_net_17             = 8'h00;
assign TX_DATA_20_const_net_17             = 8'h00;
assign TX_DATA_21_const_net_17             = 8'h00;
assign TX_DATA_22_const_net_17             = 8'h00;
assign TX_DATA_23_const_net_17             = 8'h00;
assign TX_DATA_24_const_net_17             = 8'h00;
assign TX_DATA_25_const_net_17             = 8'h00;
assign TX_DATA_26_const_net_17             = 8'h00;
assign TX_DATA_27_const_net_17             = 8'h00;
assign TX_DATA_28_const_net_17             = 8'h00;
assign TX_DATA_29_const_net_17             = 8'h00;
assign TX_DATA_30_const_net_17             = 8'h00;
assign TX_DATA_31_const_net_17             = 8'h00;
assign TX_DATA_32_const_net_17             = 8'h00;
assign TX_DATA_33_const_net_17             = 8'h00;
assign TX_DATA_34_const_net_17             = 8'h00;
assign TX_DATA_35_const_net_17             = 8'h00;
assign TX_DATA_36_const_net_17             = 8'h00;
assign TX_DATA_37_const_net_17             = 8'h00;
assign TX_DATA_38_const_net_17             = 8'h00;
assign TX_DATA_39_const_net_17             = 8'h00;
assign TX_DATA_40_const_net_17             = 8'h00;
assign TX_DATA_41_const_net_17             = 8'h00;
assign TX_DATA_42_const_net_17             = 8'h00;
assign TX_DATA_43_const_net_17             = 8'h00;
assign TX_DATA_44_const_net_17             = 8'h00;
assign TX_DATA_45_const_net_17             = 8'h00;
assign TX_DATA_46_const_net_17             = 8'h00;
assign TX_DATA_47_const_net_17             = 8'h00;
assign TX_DATA_48_const_net_17             = 8'h00;
assign TX_DATA_49_const_net_17             = 8'h00;
assign TX_DATA_50_const_net_17             = 8'h00;
assign TX_DATA_51_const_net_17             = 8'h00;
assign TX_DATA_52_const_net_17             = 8'h00;
assign TX_DATA_53_const_net_17             = 8'h00;
assign TX_DATA_54_const_net_17             = 8'h00;
assign TX_DATA_55_const_net_17             = 8'h00;
assign TX_DATA_56_const_net_17             = 8'h00;
assign TX_DATA_57_const_net_17             = 8'h00;
assign TX_DATA_58_const_net_17             = 8'h00;
assign TX_DATA_59_const_net_17             = 8'h00;
assign TX_DATA_60_const_net_17             = 8'h00;
assign TX_DATA_61_const_net_17             = 8'h00;
assign TX_DATA_62_const_net_17             = 8'h00;
assign TX_DATA_63_const_net_17             = 8'h00;
assign TX_DATA_64_const_net_17             = 8'h00;
assign TX_DATA_65_const_net_17             = 8'h00;
assign TX_DATA_66_const_net_17             = 8'h00;
assign TX_DATA_67_const_net_17             = 8'h00;
assign TX_DATA_68_const_net_17             = 8'h00;
assign TX_DATA_69_const_net_17             = 8'h00;
assign TX_DATA_70_const_net_17             = 8'h00;
assign TX_DATA_71_const_net_17             = 8'h00;
assign TX_DATA_72_const_net_17             = 8'h00;
assign TX_DATA_73_const_net_17             = 8'h00;
assign TX_DATA_74_const_net_17             = 8'h00;
assign TX_DATA_75_const_net_17             = 8'h00;
assign TX_DATA_76_const_net_17             = 8'h00;
assign TX_DATA_77_const_net_17             = 8'h00;
assign TX_DATA_78_const_net_17             = 8'h00;
assign TX_DATA_79_const_net_17             = 8'h00;
assign TX_DATA_80_const_net_17             = 8'h00;
assign TX_DATA_81_const_net_17             = 8'h00;
assign TX_DATA_82_const_net_17             = 8'h00;
assign TX_DATA_83_const_net_17             = 8'h00;
assign TX_DATA_84_const_net_17             = 8'h00;
assign TX_DATA_85_const_net_17             = 8'h00;
assign TX_DATA_86_const_net_17             = 8'h00;
assign TX_DATA_87_const_net_17             = 8'h00;
assign TX_DATA_88_const_net_17             = 8'h00;
assign TX_DATA_89_const_net_17             = 8'h00;
assign TX_DATA_90_const_net_17             = 8'h00;
assign TX_DATA_91_const_net_17             = 8'h00;
assign TX_DATA_92_const_net_17             = 8'h00;
assign TX_DATA_93_const_net_17             = 8'h00;
assign TX_DATA_94_const_net_17             = 8'h00;
assign TX_DATA_95_const_net_17             = 8'h00;
assign TX_DATA_96_const_net_17             = 8'h00;
assign TX_DATA_97_const_net_17             = 8'h00;
assign TX_DATA_98_const_net_17             = 8'h00;
assign TX_DATA_99_const_net_17             = 8'h00;
assign TX_DATA_100_const_net_17            = 8'h00;
assign TX_DATA_101_const_net_17            = 8'h00;
assign TX_DATA_102_const_net_17            = 8'h00;
assign TX_DATA_103_const_net_17            = 8'h00;
assign TX_DATA_104_const_net_17            = 8'h00;
assign TX_DATA_105_const_net_17            = 8'h00;
assign TX_DATA_106_const_net_17            = 8'h00;
assign TX_DATA_107_const_net_17            = 8'h00;
assign TX_DATA_108_const_net_17            = 8'h00;
assign TX_DATA_109_const_net_17            = 8'h00;
assign TX_DATA_110_const_net_17            = 8'h00;
assign TX_DATA_111_const_net_17            = 8'h00;
assign TX_DATA_112_const_net_17            = 8'h00;
assign TX_DATA_113_const_net_17            = 8'h00;
assign TX_DATA_114_const_net_17            = 8'h00;
assign TX_DATA_115_const_net_17            = 8'h00;
assign TX_DATA_116_const_net_17            = 8'h00;
assign TX_DATA_117_const_net_17            = 8'h00;
assign TX_DATA_118_const_net_17            = 8'h00;
assign TX_DATA_119_const_net_17            = 8'h00;
assign TX_DATA_120_const_net_17            = 8'h00;
assign TX_DATA_121_const_net_17            = 8'h00;
assign TX_DATA_122_const_net_17            = 8'h00;
assign TX_DATA_123_const_net_17            = 8'h00;
assign TX_DATA_124_const_net_17            = 8'h00;
assign TX_DATA_125_const_net_17            = 8'h00;
assign TX_DATA_126_const_net_17            = 8'h00;
assign TX_DATA_127_const_net_17            = 8'h00;
assign OE_DATA_1_const_net_16              = 4'h0;
assign OE_DATA_2_const_net_16              = 4'h0;
assign OE_DATA_3_const_net_16              = 4'h0;
assign OE_DATA_4_const_net_16              = 4'h0;
assign OE_DATA_5_const_net_16              = 4'h0;
assign OE_DATA_6_const_net_16              = 4'h0;
assign OE_DATA_7_const_net_16              = 4'h0;
assign OE_DATA_8_const_net_17              = 4'h0;
assign OE_DATA_9_const_net_17              = 4'h0;
assign OE_DATA_10_const_net_17             = 4'h0;
assign OE_DATA_11_const_net_17             = 4'h0;
assign OE_DATA_12_const_net_17             = 4'h0;
assign OE_DATA_13_const_net_17             = 4'h0;
assign OE_DATA_14_const_net_17             = 4'h0;
assign OE_DATA_15_const_net_17             = 4'h0;
assign OE_DATA_16_const_net_17             = 4'h0;
assign OE_DATA_17_const_net_17             = 4'h0;
assign OE_DATA_18_const_net_17             = 4'h0;
assign OE_DATA_19_const_net_17             = 4'h0;
assign OE_DATA_20_const_net_17             = 4'h0;
assign OE_DATA_21_const_net_17             = 4'h0;
assign OE_DATA_22_const_net_17             = 4'h0;
assign OE_DATA_23_const_net_17             = 4'h0;
assign OE_DATA_24_const_net_17             = 4'h0;
assign OE_DATA_25_const_net_17             = 4'h0;
assign OE_DATA_26_const_net_17             = 4'h0;
assign OE_DATA_27_const_net_17             = 4'h0;
assign OE_DATA_28_const_net_17             = 4'h0;
assign OE_DATA_29_const_net_17             = 4'h0;
assign OE_DATA_30_const_net_17             = 4'h0;
assign OE_DATA_31_const_net_17             = 4'h0;
assign OE_DATA_32_const_net_17             = 4'h0;
assign OE_DATA_33_const_net_17             = 4'h0;
assign OE_DATA_34_const_net_17             = 4'h0;
assign OE_DATA_35_const_net_17             = 4'h0;
assign OE_DATA_36_const_net_17             = 4'h0;
assign OE_DATA_37_const_net_17             = 4'h0;
assign OE_DATA_38_const_net_17             = 4'h0;
assign OE_DATA_39_const_net_17             = 4'h0;
assign OE_DATA_40_const_net_17             = 4'h0;
assign OE_DATA_41_const_net_17             = 4'h0;
assign OE_DATA_42_const_net_17             = 4'h0;
assign OE_DATA_43_const_net_17             = 4'h0;
assign OE_DATA_44_const_net_17             = 4'h0;
assign OE_DATA_45_const_net_17             = 4'h0;
assign OE_DATA_46_const_net_17             = 4'h0;
assign OE_DATA_47_const_net_17             = 4'h0;
assign OE_DATA_48_const_net_17             = 4'h0;
assign OE_DATA_49_const_net_17             = 4'h0;
assign OE_DATA_50_const_net_17             = 4'h0;
assign OE_DATA_51_const_net_17             = 4'h0;
assign OE_DATA_52_const_net_17             = 4'h0;
assign OE_DATA_53_const_net_17             = 4'h0;
assign OE_DATA_54_const_net_17             = 4'h0;
assign OE_DATA_55_const_net_17             = 4'h0;
assign OE_DATA_56_const_net_17             = 4'h0;
assign OE_DATA_57_const_net_17             = 4'h0;
assign OE_DATA_58_const_net_17             = 4'h0;
assign OE_DATA_59_const_net_17             = 4'h0;
assign OE_DATA_60_const_net_17             = 4'h0;
assign OE_DATA_61_const_net_17             = 4'h0;
assign OE_DATA_62_const_net_17             = 4'h0;
assign OE_DATA_63_const_net_17             = 4'h0;
assign OE_DATA_64_const_net_17             = 4'h0;
assign OE_DATA_65_const_net_17             = 4'h0;
assign OE_DATA_66_const_net_17             = 4'h0;
assign OE_DATA_67_const_net_17             = 4'h0;
assign OE_DATA_68_const_net_17             = 4'h0;
assign OE_DATA_69_const_net_17             = 4'h0;
assign OE_DATA_70_const_net_17             = 4'h0;
assign OE_DATA_71_const_net_17             = 4'h0;
assign OE_DATA_72_const_net_17             = 4'h0;
assign OE_DATA_73_const_net_17             = 4'h0;
assign OE_DATA_74_const_net_17             = 4'h0;
assign OE_DATA_75_const_net_17             = 4'h0;
assign OE_DATA_76_const_net_17             = 4'h0;
assign OE_DATA_77_const_net_17             = 4'h0;
assign OE_DATA_78_const_net_17             = 4'h0;
assign OE_DATA_79_const_net_17             = 4'h0;
assign OE_DATA_80_const_net_17             = 4'h0;
assign OE_DATA_81_const_net_17             = 4'h0;
assign OE_DATA_82_const_net_17             = 4'h0;
assign OE_DATA_83_const_net_17             = 4'h0;
assign OE_DATA_84_const_net_17             = 4'h0;
assign OE_DATA_85_const_net_17             = 4'h0;
assign OE_DATA_86_const_net_17             = 4'h0;
assign OE_DATA_87_const_net_17             = 4'h0;
assign OE_DATA_88_const_net_17             = 4'h0;
assign OE_DATA_89_const_net_17             = 4'h0;
assign OE_DATA_90_const_net_17             = 4'h0;
assign OE_DATA_91_const_net_17             = 4'h0;
assign OE_DATA_92_const_net_17             = 4'h0;
assign OE_DATA_93_const_net_17             = 4'h0;
assign OE_DATA_94_const_net_17             = 4'h0;
assign OE_DATA_95_const_net_17             = 4'h0;
assign OE_DATA_96_const_net_17             = 4'h0;
assign OE_DATA_97_const_net_17             = 4'h0;
assign OE_DATA_98_const_net_17             = 4'h0;
assign OE_DATA_99_const_net_17             = 4'h0;
assign OE_DATA_100_const_net_17            = 4'h0;
assign OE_DATA_101_const_net_17            = 4'h0;
assign OE_DATA_102_const_net_17            = 4'h0;
assign OE_DATA_103_const_net_17            = 4'h0;
assign OE_DATA_104_const_net_17            = 4'h0;
assign OE_DATA_105_const_net_17            = 4'h0;
assign OE_DATA_106_const_net_17            = 4'h0;
assign OE_DATA_107_const_net_17            = 4'h0;
assign OE_DATA_108_const_net_17            = 4'h0;
assign OE_DATA_109_const_net_17            = 4'h0;
assign OE_DATA_110_const_net_17            = 4'h0;
assign OE_DATA_111_const_net_17            = 4'h0;
assign OE_DATA_112_const_net_17            = 4'h0;
assign OE_DATA_113_const_net_17            = 4'h0;
assign OE_DATA_114_const_net_17            = 4'h0;
assign OE_DATA_115_const_net_17            = 4'h0;
assign OE_DATA_116_const_net_17            = 4'h0;
assign OE_DATA_117_const_net_17            = 4'h0;
assign OE_DATA_118_const_net_17            = 4'h0;
assign OE_DATA_119_const_net_17            = 4'h0;
assign OE_DATA_120_const_net_17            = 4'h0;
assign OE_DATA_121_const_net_17            = 4'h0;
assign OE_DATA_122_const_net_17            = 4'h0;
assign OE_DATA_123_const_net_17            = 4'h0;
assign OE_DATA_124_const_net_17            = 4'h0;
assign OE_DATA_125_const_net_17            = 4'h0;
assign OE_DATA_126_const_net_17            = 4'h0;
assign OE_DATA_127_const_net_17            = 4'h0;
assign RX_DQS_90_const_net_15              = 2'h0;
assign FIFO_WR_PTR_const_net_16            = 3'h0;
assign FIFO_RD_PTR_const_net_16            = 3'h0;
assign EYE_MONITOR_LANE_WIDTH_const_net_16 = 3'h0;
assign TX_DATA_1_const_net_14              = 2'h0;
assign TX_DATA_2_const_net_16              = 2'h0;
assign TX_DATA_3_const_net_16              = 2'h0;
assign TX_DATA_4_const_net_16              = 2'h0;
assign TX_DATA_5_const_net_16              = 2'h0;
assign TX_DATA_6_const_net_16              = 2'h0;
assign TX_DATA_7_const_net_16              = 2'h0;
assign TX_DATA_8_const_net_17              = 2'h0;
assign TX_DATA_9_const_net_17              = 2'h0;
assign TX_DATA_10_const_net_17             = 2'h0;
assign TX_DATA_11_const_net_17             = 2'h0;
assign TX_DATA_12_const_net_18             = 2'h0;
assign TX_DATA_13_const_net_18             = 2'h0;
assign TX_DATA_14_const_net_18             = 2'h0;
assign TX_DATA_15_const_net_18             = 2'h0;
assign TX_DATA_16_const_net_18             = 2'h0;
assign TX_DATA_17_const_net_18             = 2'h0;
assign TX_DATA_18_const_net_18             = 2'h0;
assign TX_DATA_19_const_net_18             = 2'h0;
assign TX_DATA_20_const_net_18             = 2'h0;
assign TX_DATA_21_const_net_18             = 2'h0;
assign TX_DATA_22_const_net_18             = 2'h0;
assign TX_DATA_23_const_net_18             = 2'h0;
assign TX_DATA_24_const_net_18             = 2'h0;
assign TX_DATA_25_const_net_18             = 2'h0;
assign TX_DATA_26_const_net_18             = 2'h0;
assign TX_DATA_27_const_net_18             = 2'h0;
assign TX_DATA_28_const_net_18             = 2'h0;
assign TX_DATA_29_const_net_18             = 2'h0;
assign TX_DATA_30_const_net_18             = 2'h0;
assign TX_DATA_31_const_net_18             = 2'h0;
assign TX_DATA_32_const_net_18             = 2'h0;
assign TX_DATA_33_const_net_18             = 2'h0;
assign TX_DATA_34_const_net_18             = 2'h0;
assign TX_DATA_35_const_net_18             = 2'h0;
assign TX_DATA_36_const_net_18             = 2'h0;
assign TX_DATA_37_const_net_18             = 2'h0;
assign TX_DATA_38_const_net_18             = 2'h0;
assign TX_DATA_39_const_net_18             = 2'h0;
assign TX_DATA_40_const_net_18             = 2'h0;
assign TX_DATA_41_const_net_18             = 2'h0;
assign TX_DATA_42_const_net_18             = 2'h0;
assign TX_DATA_43_const_net_18             = 2'h0;
assign TX_DATA_44_const_net_18             = 2'h0;
assign TX_DATA_45_const_net_18             = 2'h0;
assign TX_DATA_46_const_net_18             = 2'h0;
assign TX_DATA_47_const_net_18             = 2'h0;
assign TX_DATA_48_const_net_18             = 2'h0;
assign TX_DATA_49_const_net_18             = 2'h0;
assign TX_DATA_50_const_net_18             = 2'h0;
assign TX_DATA_51_const_net_18             = 2'h0;
assign TX_DATA_52_const_net_18             = 2'h0;
assign TX_DATA_53_const_net_18             = 2'h0;
assign TX_DATA_54_const_net_18             = 2'h0;
assign TX_DATA_55_const_net_18             = 2'h0;
assign TX_DATA_56_const_net_18             = 2'h0;
assign TX_DATA_57_const_net_18             = 2'h0;
assign TX_DATA_58_const_net_18             = 2'h0;
assign TX_DATA_59_const_net_18             = 2'h0;
assign TX_DATA_60_const_net_18             = 2'h0;
assign TX_DATA_61_const_net_18             = 2'h0;
assign TX_DATA_62_const_net_18             = 2'h0;
assign TX_DATA_63_const_net_18             = 2'h0;
assign TX_DATA_64_const_net_18             = 2'h0;
assign TX_DATA_65_const_net_18             = 2'h0;
assign TX_DATA_66_const_net_18             = 2'h0;
assign TX_DATA_67_const_net_18             = 2'h0;
assign TX_DATA_68_const_net_18             = 2'h0;
assign TX_DATA_69_const_net_18             = 2'h0;
assign TX_DATA_70_const_net_18             = 2'h0;
assign TX_DATA_71_const_net_18             = 2'h0;
assign TX_DATA_72_const_net_18             = 2'h0;
assign TX_DATA_73_const_net_18             = 2'h0;
assign TX_DATA_74_const_net_18             = 2'h0;
assign TX_DATA_75_const_net_18             = 2'h0;
assign TX_DATA_76_const_net_18             = 2'h0;
assign TX_DATA_77_const_net_18             = 2'h0;
assign TX_DATA_78_const_net_18             = 2'h0;
assign TX_DATA_79_const_net_18             = 2'h0;
assign TX_DATA_80_const_net_18             = 2'h0;
assign TX_DATA_81_const_net_18             = 2'h0;
assign TX_DATA_82_const_net_18             = 2'h0;
assign TX_DATA_83_const_net_18             = 2'h0;
assign TX_DATA_84_const_net_18             = 2'h0;
assign TX_DATA_85_const_net_18             = 2'h0;
assign TX_DATA_86_const_net_18             = 2'h0;
assign TX_DATA_87_const_net_18             = 2'h0;
assign TX_DATA_88_const_net_18             = 2'h0;
assign TX_DATA_89_const_net_18             = 2'h0;
assign TX_DATA_90_const_net_18             = 2'h0;
assign TX_DATA_91_const_net_18             = 2'h0;
assign TX_DATA_92_const_net_18             = 2'h0;
assign TX_DATA_93_const_net_18             = 2'h0;
assign TX_DATA_94_const_net_18             = 2'h0;
assign TX_DATA_95_const_net_18             = 2'h0;
assign TX_DATA_96_const_net_18             = 2'h0;
assign TX_DATA_97_const_net_18             = 2'h0;
assign TX_DATA_98_const_net_18             = 2'h0;
assign TX_DATA_99_const_net_18             = 2'h0;
assign TX_DATA_100_const_net_18            = 2'h0;
assign TX_DATA_101_const_net_18            = 2'h0;
assign TX_DATA_102_const_net_18            = 2'h0;
assign TX_DATA_103_const_net_18            = 2'h0;
assign TX_DATA_104_const_net_18            = 2'h0;
assign TX_DATA_105_const_net_18            = 2'h0;
assign TX_DATA_106_const_net_18            = 2'h0;
assign TX_DATA_107_const_net_18            = 2'h0;
assign TX_DATA_108_const_net_18            = 2'h0;
assign TX_DATA_109_const_net_18            = 2'h0;
assign TX_DATA_110_const_net_18            = 2'h0;
assign TX_DATA_111_const_net_18            = 2'h0;
assign TX_DATA_112_const_net_18            = 2'h0;
assign TX_DATA_113_const_net_18            = 2'h0;
assign TX_DATA_114_const_net_18            = 2'h0;
assign TX_DATA_115_const_net_18            = 2'h0;
assign TX_DATA_116_const_net_18            = 2'h0;
assign TX_DATA_117_const_net_18            = 2'h0;
assign TX_DATA_118_const_net_18            = 2'h0;
assign TX_DATA_119_const_net_18            = 2'h0;
assign TX_DATA_120_const_net_18            = 2'h0;
assign TX_DATA_121_const_net_18            = 2'h0;
assign TX_DATA_122_const_net_18            = 2'h0;
assign TX_DATA_123_const_net_18            = 2'h0;
assign TX_DATA_124_const_net_18            = 2'h0;
assign TX_DATA_125_const_net_18            = 2'h0;
assign TX_DATA_126_const_net_18            = 2'h0;
assign TX_DATA_127_const_net_18            = 2'h0;
assign OE_DATA_1_const_net_17              = 2'h0;
assign OE_DATA_2_const_net_17              = 2'h0;
assign OE_DATA_3_const_net_17              = 2'h0;
assign OE_DATA_4_const_net_17              = 2'h0;
assign OE_DATA_5_const_net_17              = 2'h0;
assign OE_DATA_6_const_net_17              = 2'h0;
assign OE_DATA_7_const_net_17              = 2'h0;
assign OE_DATA_8_const_net_18              = 2'h0;
assign OE_DATA_9_const_net_18              = 2'h0;
assign OE_DATA_10_const_net_18             = 2'h0;
assign OE_DATA_11_const_net_18             = 2'h0;
assign OE_DATA_12_const_net_18             = 2'h0;
assign OE_DATA_13_const_net_18             = 2'h0;
assign OE_DATA_14_const_net_18             = 2'h0;
assign OE_DATA_15_const_net_18             = 2'h0;
assign OE_DATA_16_const_net_18             = 2'h0;
assign OE_DATA_17_const_net_18             = 2'h0;
assign OE_DATA_18_const_net_18             = 2'h0;
assign OE_DATA_19_const_net_18             = 2'h0;
assign OE_DATA_20_const_net_18             = 2'h0;
assign OE_DATA_21_const_net_18             = 2'h0;
assign OE_DATA_22_const_net_18             = 2'h0;
assign OE_DATA_23_const_net_18             = 2'h0;
assign OE_DATA_24_const_net_18             = 2'h0;
assign OE_DATA_25_const_net_18             = 2'h0;
assign OE_DATA_26_const_net_18             = 2'h0;
assign OE_DATA_27_const_net_18             = 2'h0;
assign OE_DATA_28_const_net_18             = 2'h0;
assign OE_DATA_29_const_net_18             = 2'h0;
assign OE_DATA_30_const_net_18             = 2'h0;
assign OE_DATA_31_const_net_18             = 2'h0;
assign OE_DATA_32_const_net_18             = 2'h0;
assign OE_DATA_33_const_net_18             = 2'h0;
assign OE_DATA_34_const_net_18             = 2'h0;
assign OE_DATA_35_const_net_18             = 2'h0;
assign OE_DATA_36_const_net_18             = 2'h0;
assign OE_DATA_37_const_net_18             = 2'h0;
assign OE_DATA_38_const_net_18             = 2'h0;
assign OE_DATA_39_const_net_18             = 2'h0;
assign OE_DATA_40_const_net_18             = 2'h0;
assign OE_DATA_41_const_net_18             = 2'h0;
assign OE_DATA_42_const_net_18             = 2'h0;
assign OE_DATA_43_const_net_18             = 2'h0;
assign OE_DATA_44_const_net_18             = 2'h0;
assign OE_DATA_45_const_net_18             = 2'h0;
assign OE_DATA_46_const_net_18             = 2'h0;
assign OE_DATA_47_const_net_18             = 2'h0;
assign OE_DATA_48_const_net_18             = 2'h0;
assign OE_DATA_49_const_net_18             = 2'h0;
assign OE_DATA_50_const_net_18             = 2'h0;
assign OE_DATA_51_const_net_18             = 2'h0;
assign OE_DATA_52_const_net_18             = 2'h0;
assign OE_DATA_53_const_net_18             = 2'h0;
assign OE_DATA_54_const_net_18             = 2'h0;
assign OE_DATA_55_const_net_18             = 2'h0;
assign OE_DATA_56_const_net_18             = 2'h0;
assign OE_DATA_57_const_net_18             = 2'h0;
assign OE_DATA_58_const_net_18             = 2'h0;
assign OE_DATA_59_const_net_18             = 2'h0;
assign OE_DATA_60_const_net_18             = 2'h0;
assign OE_DATA_61_const_net_18             = 2'h0;
assign OE_DATA_62_const_net_18             = 2'h0;
assign OE_DATA_63_const_net_18             = 2'h0;
assign OE_DATA_64_const_net_18             = 2'h0;
assign OE_DATA_65_const_net_18             = 2'h0;
assign OE_DATA_66_const_net_18             = 2'h0;
assign OE_DATA_67_const_net_18             = 2'h0;
assign OE_DATA_68_const_net_18             = 2'h0;
assign OE_DATA_69_const_net_18             = 2'h0;
assign OE_DATA_70_const_net_18             = 2'h0;
assign OE_DATA_71_const_net_18             = 2'h0;
assign OE_DATA_72_const_net_18             = 2'h0;
assign OE_DATA_73_const_net_18             = 2'h0;
assign OE_DATA_74_const_net_18             = 2'h0;
assign OE_DATA_75_const_net_18             = 2'h0;
assign OE_DATA_76_const_net_18             = 2'h0;
assign OE_DATA_77_const_net_18             = 2'h0;
assign OE_DATA_78_const_net_18             = 2'h0;
assign OE_DATA_79_const_net_18             = 2'h0;
assign OE_DATA_80_const_net_18             = 2'h0;
assign OE_DATA_81_const_net_18             = 2'h0;
assign OE_DATA_82_const_net_18             = 2'h0;
assign OE_DATA_83_const_net_18             = 2'h0;
assign OE_DATA_84_const_net_18             = 2'h0;
assign OE_DATA_85_const_net_18             = 2'h0;
assign OE_DATA_86_const_net_18             = 2'h0;
assign OE_DATA_87_const_net_18             = 2'h0;
assign OE_DATA_88_const_net_18             = 2'h0;
assign OE_DATA_89_const_net_18             = 2'h0;
assign OE_DATA_90_const_net_18             = 2'h0;
assign OE_DATA_91_const_net_18             = 2'h0;
assign OE_DATA_92_const_net_18             = 2'h0;
assign OE_DATA_93_const_net_18             = 2'h0;
assign OE_DATA_94_const_net_18             = 2'h0;
assign OE_DATA_95_const_net_18             = 2'h0;
assign OE_DATA_96_const_net_18             = 2'h0;
assign OE_DATA_97_const_net_18             = 2'h0;
assign OE_DATA_98_const_net_18             = 2'h0;
assign OE_DATA_99_const_net_18             = 2'h0;
assign OE_DATA_100_const_net_18            = 2'h0;
assign OE_DATA_101_const_net_18            = 2'h0;
assign OE_DATA_102_const_net_18            = 2'h0;
assign OE_DATA_103_const_net_18            = 2'h0;
assign OE_DATA_104_const_net_18            = 2'h0;
assign OE_DATA_105_const_net_18            = 2'h0;
assign OE_DATA_106_const_net_18            = 2'h0;
assign OE_DATA_107_const_net_18            = 2'h0;
assign OE_DATA_108_const_net_18            = 2'h0;
assign OE_DATA_109_const_net_18            = 2'h0;
assign OE_DATA_110_const_net_18            = 2'h0;
assign OE_DATA_111_const_net_18            = 2'h0;
assign OE_DATA_112_const_net_18            = 2'h0;
assign OE_DATA_113_const_net_18            = 2'h0;
assign OE_DATA_114_const_net_18            = 2'h0;
assign OE_DATA_115_const_net_18            = 2'h0;
assign OE_DATA_116_const_net_18            = 2'h0;
assign OE_DATA_117_const_net_18            = 2'h0;
assign OE_DATA_118_const_net_18            = 2'h0;
assign OE_DATA_119_const_net_18            = 2'h0;
assign OE_DATA_120_const_net_18            = 2'h0;
assign OE_DATA_121_const_net_18            = 2'h0;
assign OE_DATA_122_const_net_18            = 2'h0;
assign OE_DATA_123_const_net_18            = 2'h0;
assign OE_DATA_124_const_net_18            = 2'h0;
assign OE_DATA_125_const_net_18            = 2'h0;
assign OE_DATA_126_const_net_18            = 2'h0;
assign OE_DATA_127_const_net_18            = 2'h0;
assign RX_DQS_90_const_net_16              = 2'h0;
assign EYE_MONITOR_LANE_WIDTH_const_net_17 = 3'h0;
assign TX_DATA_1_const_net_15              = 8'h00;
assign TX_DATA_2_const_net_17              = 8'h00;
assign TX_DATA_3_const_net_17              = 8'h00;
assign TX_DATA_4_const_net_17              = 8'h00;
assign TX_DATA_5_const_net_17              = 8'h00;
assign TX_DATA_6_const_net_17              = 8'h00;
assign TX_DATA_7_const_net_17              = 8'h00;
assign TX_DATA_8_const_net_18              = 8'h00;
assign TX_DATA_9_const_net_18              = 8'h00;
assign TX_DATA_10_const_net_18             = 8'h00;
assign TX_DATA_11_const_net_18             = 8'h00;
assign TX_DATA_12_const_net_19             = 8'h00;
assign TX_DATA_13_const_net_19             = 8'h00;
assign TX_DATA_14_const_net_19             = 8'h00;
assign TX_DATA_15_const_net_19             = 8'h00;
assign TX_DATA_16_const_net_19             = 8'h00;
assign TX_DATA_17_const_net_19             = 8'h00;
assign TX_DATA_18_const_net_19             = 8'h00;
assign TX_DATA_19_const_net_19             = 8'h00;
assign TX_DATA_20_const_net_19             = 8'h00;
assign TX_DATA_21_const_net_19             = 8'h00;
assign TX_DATA_22_const_net_19             = 8'h00;
assign TX_DATA_23_const_net_19             = 8'h00;
assign TX_DATA_24_const_net_19             = 8'h00;
assign TX_DATA_25_const_net_19             = 8'h00;
assign TX_DATA_26_const_net_19             = 8'h00;
assign TX_DATA_27_const_net_19             = 8'h00;
assign TX_DATA_28_const_net_19             = 8'h00;
assign TX_DATA_29_const_net_19             = 8'h00;
assign TX_DATA_30_const_net_19             = 8'h00;
assign TX_DATA_31_const_net_19             = 8'h00;
assign TX_DATA_32_const_net_19             = 8'h00;
assign TX_DATA_33_const_net_19             = 8'h00;
assign TX_DATA_34_const_net_19             = 8'h00;
assign TX_DATA_35_const_net_19             = 8'h00;
assign TX_DATA_36_const_net_19             = 8'h00;
assign TX_DATA_37_const_net_19             = 8'h00;
assign TX_DATA_38_const_net_19             = 8'h00;
assign TX_DATA_39_const_net_19             = 8'h00;
assign TX_DATA_40_const_net_19             = 8'h00;
assign TX_DATA_41_const_net_19             = 8'h00;
assign TX_DATA_42_const_net_19             = 8'h00;
assign TX_DATA_43_const_net_19             = 8'h00;
assign TX_DATA_44_const_net_19             = 8'h00;
assign TX_DATA_45_const_net_19             = 8'h00;
assign TX_DATA_46_const_net_19             = 8'h00;
assign TX_DATA_47_const_net_19             = 8'h00;
assign TX_DATA_48_const_net_19             = 8'h00;
assign TX_DATA_49_const_net_19             = 8'h00;
assign TX_DATA_50_const_net_19             = 8'h00;
assign TX_DATA_51_const_net_19             = 8'h00;
assign TX_DATA_52_const_net_19             = 8'h00;
assign TX_DATA_53_const_net_19             = 8'h00;
assign TX_DATA_54_const_net_19             = 8'h00;
assign TX_DATA_55_const_net_19             = 8'h00;
assign TX_DATA_56_const_net_19             = 8'h00;
assign TX_DATA_57_const_net_19             = 8'h00;
assign TX_DATA_58_const_net_19             = 8'h00;
assign TX_DATA_59_const_net_19             = 8'h00;
assign TX_DATA_60_const_net_19             = 8'h00;
assign TX_DATA_61_const_net_19             = 8'h00;
assign TX_DATA_62_const_net_19             = 8'h00;
assign TX_DATA_63_const_net_19             = 8'h00;
assign TX_DATA_64_const_net_19             = 8'h00;
assign TX_DATA_65_const_net_19             = 8'h00;
assign TX_DATA_66_const_net_19             = 8'h00;
assign TX_DATA_67_const_net_19             = 8'h00;
assign TX_DATA_68_const_net_19             = 8'h00;
assign TX_DATA_69_const_net_19             = 8'h00;
assign TX_DATA_70_const_net_19             = 8'h00;
assign TX_DATA_71_const_net_19             = 8'h00;
assign TX_DATA_72_const_net_19             = 8'h00;
assign TX_DATA_73_const_net_19             = 8'h00;
assign TX_DATA_74_const_net_19             = 8'h00;
assign TX_DATA_75_const_net_19             = 8'h00;
assign TX_DATA_76_const_net_19             = 8'h00;
assign TX_DATA_77_const_net_19             = 8'h00;
assign TX_DATA_78_const_net_19             = 8'h00;
assign TX_DATA_79_const_net_19             = 8'h00;
assign TX_DATA_80_const_net_19             = 8'h00;
assign TX_DATA_81_const_net_19             = 8'h00;
assign TX_DATA_82_const_net_19             = 8'h00;
assign TX_DATA_83_const_net_19             = 8'h00;
assign TX_DATA_84_const_net_19             = 8'h00;
assign TX_DATA_85_const_net_19             = 8'h00;
assign TX_DATA_86_const_net_19             = 8'h00;
assign TX_DATA_87_const_net_19             = 8'h00;
assign TX_DATA_88_const_net_19             = 8'h00;
assign TX_DATA_89_const_net_19             = 8'h00;
assign TX_DATA_90_const_net_19             = 8'h00;
assign TX_DATA_91_const_net_19             = 8'h00;
assign TX_DATA_92_const_net_19             = 8'h00;
assign TX_DATA_93_const_net_19             = 8'h00;
assign TX_DATA_94_const_net_19             = 8'h00;
assign TX_DATA_95_const_net_19             = 8'h00;
assign TX_DATA_96_const_net_19             = 8'h00;
assign TX_DATA_97_const_net_19             = 8'h00;
assign TX_DATA_98_const_net_19             = 8'h00;
assign TX_DATA_99_const_net_19             = 8'h00;
assign TX_DATA_100_const_net_19            = 8'h00;
assign TX_DATA_101_const_net_19            = 8'h00;
assign TX_DATA_102_const_net_19            = 8'h00;
assign TX_DATA_103_const_net_19            = 8'h00;
assign TX_DATA_104_const_net_19            = 8'h00;
assign TX_DATA_105_const_net_19            = 8'h00;
assign TX_DATA_106_const_net_19            = 8'h00;
assign TX_DATA_107_const_net_19            = 8'h00;
assign TX_DATA_108_const_net_19            = 8'h00;
assign TX_DATA_109_const_net_19            = 8'h00;
assign TX_DATA_110_const_net_19            = 8'h00;
assign TX_DATA_111_const_net_19            = 8'h00;
assign TX_DATA_112_const_net_19            = 8'h00;
assign TX_DATA_113_const_net_19            = 8'h00;
assign TX_DATA_114_const_net_19            = 8'h00;
assign TX_DATA_115_const_net_19            = 8'h00;
assign TX_DATA_116_const_net_19            = 8'h00;
assign TX_DATA_117_const_net_19            = 8'h00;
assign TX_DATA_118_const_net_19            = 8'h00;
assign TX_DATA_119_const_net_19            = 8'h00;
assign TX_DATA_120_const_net_19            = 8'h00;
assign TX_DATA_121_const_net_19            = 8'h00;
assign TX_DATA_122_const_net_19            = 8'h00;
assign TX_DATA_123_const_net_19            = 8'h00;
assign TX_DATA_124_const_net_19            = 8'h00;
assign TX_DATA_125_const_net_19            = 8'h00;
assign TX_DATA_126_const_net_19            = 8'h00;
assign TX_DATA_127_const_net_19            = 8'h00;
assign OE_DATA_1_const_net_18              = 4'h0;
assign OE_DATA_2_const_net_18              = 4'h0;
assign OE_DATA_3_const_net_18              = 4'h0;
assign OE_DATA_4_const_net_18              = 4'h0;
assign OE_DATA_5_const_net_18              = 4'h0;
assign OE_DATA_6_const_net_18              = 4'h0;
assign OE_DATA_7_const_net_18              = 4'h0;
assign OE_DATA_8_const_net_19              = 4'h0;
assign OE_DATA_9_const_net_19              = 4'h0;
assign OE_DATA_10_const_net_19             = 4'h0;
assign OE_DATA_11_const_net_19             = 4'h0;
assign OE_DATA_12_const_net_19             = 4'h0;
assign OE_DATA_13_const_net_19             = 4'h0;
assign OE_DATA_14_const_net_19             = 4'h0;
assign OE_DATA_15_const_net_19             = 4'h0;
assign OE_DATA_16_const_net_19             = 4'h0;
assign OE_DATA_17_const_net_19             = 4'h0;
assign OE_DATA_18_const_net_19             = 4'h0;
assign OE_DATA_19_const_net_19             = 4'h0;
assign OE_DATA_20_const_net_19             = 4'h0;
assign OE_DATA_21_const_net_19             = 4'h0;
assign OE_DATA_22_const_net_19             = 4'h0;
assign OE_DATA_23_const_net_19             = 4'h0;
assign OE_DATA_24_const_net_19             = 4'h0;
assign OE_DATA_25_const_net_19             = 4'h0;
assign OE_DATA_26_const_net_19             = 4'h0;
assign OE_DATA_27_const_net_19             = 4'h0;
assign OE_DATA_28_const_net_19             = 4'h0;
assign OE_DATA_29_const_net_19             = 4'h0;
assign OE_DATA_30_const_net_19             = 4'h0;
assign OE_DATA_31_const_net_19             = 4'h0;
assign OE_DATA_32_const_net_19             = 4'h0;
assign OE_DATA_33_const_net_19             = 4'h0;
assign OE_DATA_34_const_net_19             = 4'h0;
assign OE_DATA_35_const_net_19             = 4'h0;
assign OE_DATA_36_const_net_19             = 4'h0;
assign OE_DATA_37_const_net_19             = 4'h0;
assign OE_DATA_38_const_net_19             = 4'h0;
assign OE_DATA_39_const_net_19             = 4'h0;
assign OE_DATA_40_const_net_19             = 4'h0;
assign OE_DATA_41_const_net_19             = 4'h0;
assign OE_DATA_42_const_net_19             = 4'h0;
assign OE_DATA_43_const_net_19             = 4'h0;
assign OE_DATA_44_const_net_19             = 4'h0;
assign OE_DATA_45_const_net_19             = 4'h0;
assign OE_DATA_46_const_net_19             = 4'h0;
assign OE_DATA_47_const_net_19             = 4'h0;
assign OE_DATA_48_const_net_19             = 4'h0;
assign OE_DATA_49_const_net_19             = 4'h0;
assign OE_DATA_50_const_net_19             = 4'h0;
assign OE_DATA_51_const_net_19             = 4'h0;
assign OE_DATA_52_const_net_19             = 4'h0;
assign OE_DATA_53_const_net_19             = 4'h0;
assign OE_DATA_54_const_net_19             = 4'h0;
assign OE_DATA_55_const_net_19             = 4'h0;
assign OE_DATA_56_const_net_19             = 4'h0;
assign OE_DATA_57_const_net_19             = 4'h0;
assign OE_DATA_58_const_net_19             = 4'h0;
assign OE_DATA_59_const_net_19             = 4'h0;
assign OE_DATA_60_const_net_19             = 4'h0;
assign OE_DATA_61_const_net_19             = 4'h0;
assign OE_DATA_62_const_net_19             = 4'h0;
assign OE_DATA_63_const_net_19             = 4'h0;
assign OE_DATA_64_const_net_19             = 4'h0;
assign OE_DATA_65_const_net_19             = 4'h0;
assign OE_DATA_66_const_net_19             = 4'h0;
assign OE_DATA_67_const_net_19             = 4'h0;
assign OE_DATA_68_const_net_19             = 4'h0;
assign OE_DATA_69_const_net_19             = 4'h0;
assign OE_DATA_70_const_net_19             = 4'h0;
assign OE_DATA_71_const_net_19             = 4'h0;
assign OE_DATA_72_const_net_19             = 4'h0;
assign OE_DATA_73_const_net_19             = 4'h0;
assign OE_DATA_74_const_net_19             = 4'h0;
assign OE_DATA_75_const_net_19             = 4'h0;
assign OE_DATA_76_const_net_19             = 4'h0;
assign OE_DATA_77_const_net_19             = 4'h0;
assign OE_DATA_78_const_net_19             = 4'h0;
assign OE_DATA_79_const_net_19             = 4'h0;
assign OE_DATA_80_const_net_19             = 4'h0;
assign OE_DATA_81_const_net_19             = 4'h0;
assign OE_DATA_82_const_net_19             = 4'h0;
assign OE_DATA_83_const_net_19             = 4'h0;
assign OE_DATA_84_const_net_19             = 4'h0;
assign OE_DATA_85_const_net_19             = 4'h0;
assign OE_DATA_86_const_net_19             = 4'h0;
assign OE_DATA_87_const_net_19             = 4'h0;
assign OE_DATA_88_const_net_19             = 4'h0;
assign OE_DATA_89_const_net_19             = 4'h0;
assign OE_DATA_90_const_net_19             = 4'h0;
assign OE_DATA_91_const_net_19             = 4'h0;
assign OE_DATA_92_const_net_19             = 4'h0;
assign OE_DATA_93_const_net_19             = 4'h0;
assign OE_DATA_94_const_net_19             = 4'h0;
assign OE_DATA_95_const_net_19             = 4'h0;
assign OE_DATA_96_const_net_19             = 4'h0;
assign OE_DATA_97_const_net_19             = 4'h0;
assign OE_DATA_98_const_net_19             = 4'h0;
assign OE_DATA_99_const_net_19             = 4'h0;
assign OE_DATA_100_const_net_19            = 4'h0;
assign OE_DATA_101_const_net_19            = 4'h0;
assign OE_DATA_102_const_net_19            = 4'h0;
assign OE_DATA_103_const_net_19            = 4'h0;
assign OE_DATA_104_const_net_19            = 4'h0;
assign OE_DATA_105_const_net_19            = 4'h0;
assign OE_DATA_106_const_net_19            = 4'h0;
assign OE_DATA_107_const_net_19            = 4'h0;
assign OE_DATA_108_const_net_19            = 4'h0;
assign OE_DATA_109_const_net_19            = 4'h0;
assign OE_DATA_110_const_net_19            = 4'h0;
assign OE_DATA_111_const_net_19            = 4'h0;
assign OE_DATA_112_const_net_19            = 4'h0;
assign OE_DATA_113_const_net_19            = 4'h0;
assign OE_DATA_114_const_net_19            = 4'h0;
assign OE_DATA_115_const_net_19            = 4'h0;
assign OE_DATA_116_const_net_19            = 4'h0;
assign OE_DATA_117_const_net_19            = 4'h0;
assign OE_DATA_118_const_net_19            = 4'h0;
assign OE_DATA_119_const_net_19            = 4'h0;
assign OE_DATA_120_const_net_19            = 4'h0;
assign OE_DATA_121_const_net_19            = 4'h0;
assign OE_DATA_122_const_net_19            = 4'h0;
assign OE_DATA_123_const_net_19            = 4'h0;
assign OE_DATA_124_const_net_19            = 4'h0;
assign OE_DATA_125_const_net_19            = 4'h0;
assign OE_DATA_126_const_net_19            = 4'h0;
assign OE_DATA_127_const_net_19            = 4'h0;
assign CDR_CLK_B_SEL_const_net_1           = 11'h000;
assign FIFO_WR_PTR_const_net_17            = 3'h0;
assign FIFO_RD_PTR_const_net_17            = 3'h0;
assign EYE_MONITOR_LANE_WIDTH_const_net_18 = 3'h0;
assign TX_DATA_1_const_net_16              = 8'h00;
assign TX_DATA_2_const_net_18              = 8'h00;
assign TX_DATA_3_const_net_18              = 8'h00;
assign TX_DATA_4_const_net_18              = 8'h00;
assign TX_DATA_5_const_net_18              = 8'h00;
assign TX_DATA_6_const_net_18              = 8'h00;
assign TX_DATA_7_const_net_18              = 8'h00;
assign TX_DATA_8_const_net_19              = 8'h00;
assign TX_DATA_9_const_net_19              = 8'h00;
assign TX_DATA_10_const_net_19             = 8'h00;
assign TX_DATA_11_const_net_19             = 8'h00;
assign TX_DATA_12_const_net_20             = 8'h00;
assign TX_DATA_13_const_net_20             = 8'h00;
assign TX_DATA_14_const_net_20             = 8'h00;
assign TX_DATA_15_const_net_20             = 8'h00;
assign TX_DATA_16_const_net_20             = 8'h00;
assign TX_DATA_17_const_net_20             = 8'h00;
assign TX_DATA_18_const_net_20             = 8'h00;
assign TX_DATA_19_const_net_20             = 8'h00;
assign TX_DATA_20_const_net_20             = 8'h00;
assign TX_DATA_21_const_net_20             = 8'h00;
assign TX_DATA_22_const_net_20             = 8'h00;
assign TX_DATA_23_const_net_20             = 8'h00;
assign TX_DATA_24_const_net_20             = 8'h00;
assign TX_DATA_25_const_net_20             = 8'h00;
assign TX_DATA_26_const_net_20             = 8'h00;
assign TX_DATA_27_const_net_20             = 8'h00;
assign TX_DATA_28_const_net_20             = 8'h00;
assign TX_DATA_29_const_net_20             = 8'h00;
assign TX_DATA_30_const_net_20             = 8'h00;
assign TX_DATA_31_const_net_20             = 8'h00;
assign TX_DATA_32_const_net_20             = 8'h00;
assign TX_DATA_33_const_net_20             = 8'h00;
assign TX_DATA_34_const_net_20             = 8'h00;
assign TX_DATA_35_const_net_20             = 8'h00;
assign TX_DATA_36_const_net_20             = 8'h00;
assign TX_DATA_37_const_net_20             = 8'h00;
assign TX_DATA_38_const_net_20             = 8'h00;
assign TX_DATA_39_const_net_20             = 8'h00;
assign TX_DATA_40_const_net_20             = 8'h00;
assign TX_DATA_41_const_net_20             = 8'h00;
assign TX_DATA_42_const_net_20             = 8'h00;
assign TX_DATA_43_const_net_20             = 8'h00;
assign TX_DATA_44_const_net_20             = 8'h00;
assign TX_DATA_45_const_net_20             = 8'h00;
assign TX_DATA_46_const_net_20             = 8'h00;
assign TX_DATA_47_const_net_20             = 8'h00;
assign TX_DATA_48_const_net_20             = 8'h00;
assign TX_DATA_49_const_net_20             = 8'h00;
assign TX_DATA_50_const_net_20             = 8'h00;
assign TX_DATA_51_const_net_20             = 8'h00;
assign TX_DATA_52_const_net_20             = 8'h00;
assign TX_DATA_53_const_net_20             = 8'h00;
assign TX_DATA_54_const_net_20             = 8'h00;
assign TX_DATA_55_const_net_20             = 8'h00;
assign TX_DATA_56_const_net_20             = 8'h00;
assign TX_DATA_57_const_net_20             = 8'h00;
assign TX_DATA_58_const_net_20             = 8'h00;
assign TX_DATA_59_const_net_20             = 8'h00;
assign TX_DATA_60_const_net_20             = 8'h00;
assign TX_DATA_61_const_net_20             = 8'h00;
assign TX_DATA_62_const_net_20             = 8'h00;
assign TX_DATA_63_const_net_20             = 8'h00;
assign TX_DATA_64_const_net_20             = 8'h00;
assign TX_DATA_65_const_net_20             = 8'h00;
assign TX_DATA_66_const_net_20             = 8'h00;
assign TX_DATA_67_const_net_20             = 8'h00;
assign TX_DATA_68_const_net_20             = 8'h00;
assign TX_DATA_69_const_net_20             = 8'h00;
assign TX_DATA_70_const_net_20             = 8'h00;
assign TX_DATA_71_const_net_20             = 8'h00;
assign TX_DATA_72_const_net_20             = 8'h00;
assign TX_DATA_73_const_net_20             = 8'h00;
assign TX_DATA_74_const_net_20             = 8'h00;
assign TX_DATA_75_const_net_20             = 8'h00;
assign TX_DATA_76_const_net_20             = 8'h00;
assign TX_DATA_77_const_net_20             = 8'h00;
assign TX_DATA_78_const_net_20             = 8'h00;
assign TX_DATA_79_const_net_20             = 8'h00;
assign TX_DATA_80_const_net_20             = 8'h00;
assign TX_DATA_81_const_net_20             = 8'h00;
assign TX_DATA_82_const_net_20             = 8'h00;
assign TX_DATA_83_const_net_20             = 8'h00;
assign TX_DATA_84_const_net_20             = 8'h00;
assign TX_DATA_85_const_net_20             = 8'h00;
assign TX_DATA_86_const_net_20             = 8'h00;
assign TX_DATA_87_const_net_20             = 8'h00;
assign TX_DATA_88_const_net_20             = 8'h00;
assign TX_DATA_89_const_net_20             = 8'h00;
assign TX_DATA_90_const_net_20             = 8'h00;
assign TX_DATA_91_const_net_20             = 8'h00;
assign TX_DATA_92_const_net_20             = 8'h00;
assign TX_DATA_93_const_net_20             = 8'h00;
assign TX_DATA_94_const_net_20             = 8'h00;
assign TX_DATA_95_const_net_20             = 8'h00;
assign TX_DATA_96_const_net_20             = 8'h00;
assign TX_DATA_97_const_net_20             = 8'h00;
assign TX_DATA_98_const_net_20             = 8'h00;
assign TX_DATA_99_const_net_20             = 8'h00;
assign TX_DATA_100_const_net_20            = 8'h00;
assign TX_DATA_101_const_net_20            = 8'h00;
assign TX_DATA_102_const_net_20            = 8'h00;
assign TX_DATA_103_const_net_20            = 8'h00;
assign TX_DATA_104_const_net_20            = 8'h00;
assign TX_DATA_105_const_net_20            = 8'h00;
assign TX_DATA_106_const_net_20            = 8'h00;
assign TX_DATA_107_const_net_20            = 8'h00;
assign TX_DATA_108_const_net_20            = 8'h00;
assign TX_DATA_109_const_net_20            = 8'h00;
assign TX_DATA_110_const_net_20            = 8'h00;
assign TX_DATA_111_const_net_20            = 8'h00;
assign TX_DATA_112_const_net_20            = 8'h00;
assign TX_DATA_113_const_net_20            = 8'h00;
assign TX_DATA_114_const_net_20            = 8'h00;
assign TX_DATA_115_const_net_20            = 8'h00;
assign TX_DATA_116_const_net_20            = 8'h00;
assign TX_DATA_117_const_net_20            = 8'h00;
assign TX_DATA_118_const_net_20            = 8'h00;
assign TX_DATA_119_const_net_20            = 8'h00;
assign TX_DATA_120_const_net_20            = 8'h00;
assign TX_DATA_121_const_net_20            = 8'h00;
assign TX_DATA_122_const_net_20            = 8'h00;
assign TX_DATA_123_const_net_20            = 8'h00;
assign TX_DATA_124_const_net_20            = 8'h00;
assign TX_DATA_125_const_net_20            = 8'h00;
assign TX_DATA_126_const_net_20            = 8'h00;
assign TX_DATA_127_const_net_20            = 8'h00;
assign OE_DATA_1_const_net_19              = 4'h0;
assign OE_DATA_2_const_net_19              = 4'h0;
assign OE_DATA_3_const_net_19              = 4'h0;
assign OE_DATA_4_const_net_19              = 4'h0;
assign OE_DATA_5_const_net_19              = 4'h0;
assign OE_DATA_6_const_net_19              = 4'h0;
assign OE_DATA_7_const_net_19              = 4'h0;
assign OE_DATA_8_const_net_20              = 4'h0;
assign OE_DATA_9_const_net_20              = 4'h0;
assign OE_DATA_10_const_net_20             = 4'h0;
assign OE_DATA_11_const_net_20             = 4'h0;
assign OE_DATA_12_const_net_20             = 4'h0;
assign OE_DATA_13_const_net_20             = 4'h0;
assign OE_DATA_14_const_net_20             = 4'h0;
assign OE_DATA_15_const_net_20             = 4'h0;
assign OE_DATA_16_const_net_20             = 4'h0;
assign OE_DATA_17_const_net_20             = 4'h0;
assign OE_DATA_18_const_net_20             = 4'h0;
assign OE_DATA_19_const_net_20             = 4'h0;
assign OE_DATA_20_const_net_20             = 4'h0;
assign OE_DATA_21_const_net_20             = 4'h0;
assign OE_DATA_22_const_net_20             = 4'h0;
assign OE_DATA_23_const_net_20             = 4'h0;
assign OE_DATA_24_const_net_20             = 4'h0;
assign OE_DATA_25_const_net_20             = 4'h0;
assign OE_DATA_26_const_net_20             = 4'h0;
assign OE_DATA_27_const_net_20             = 4'h0;
assign OE_DATA_28_const_net_20             = 4'h0;
assign OE_DATA_29_const_net_20             = 4'h0;
assign OE_DATA_30_const_net_20             = 4'h0;
assign OE_DATA_31_const_net_20             = 4'h0;
assign OE_DATA_32_const_net_20             = 4'h0;
assign OE_DATA_33_const_net_20             = 4'h0;
assign OE_DATA_34_const_net_20             = 4'h0;
assign OE_DATA_35_const_net_20             = 4'h0;
assign OE_DATA_36_const_net_20             = 4'h0;
assign OE_DATA_37_const_net_20             = 4'h0;
assign OE_DATA_38_const_net_20             = 4'h0;
assign OE_DATA_39_const_net_20             = 4'h0;
assign OE_DATA_40_const_net_20             = 4'h0;
assign OE_DATA_41_const_net_20             = 4'h0;
assign OE_DATA_42_const_net_20             = 4'h0;
assign OE_DATA_43_const_net_20             = 4'h0;
assign OE_DATA_44_const_net_20             = 4'h0;
assign OE_DATA_45_const_net_20             = 4'h0;
assign OE_DATA_46_const_net_20             = 4'h0;
assign OE_DATA_47_const_net_20             = 4'h0;
assign OE_DATA_48_const_net_20             = 4'h0;
assign OE_DATA_49_const_net_20             = 4'h0;
assign OE_DATA_50_const_net_20             = 4'h0;
assign OE_DATA_51_const_net_20             = 4'h0;
assign OE_DATA_52_const_net_20             = 4'h0;
assign OE_DATA_53_const_net_20             = 4'h0;
assign OE_DATA_54_const_net_20             = 4'h0;
assign OE_DATA_55_const_net_20             = 4'h0;
assign OE_DATA_56_const_net_20             = 4'h0;
assign OE_DATA_57_const_net_20             = 4'h0;
assign OE_DATA_58_const_net_20             = 4'h0;
assign OE_DATA_59_const_net_20             = 4'h0;
assign OE_DATA_60_const_net_20             = 4'h0;
assign OE_DATA_61_const_net_20             = 4'h0;
assign OE_DATA_62_const_net_20             = 4'h0;
assign OE_DATA_63_const_net_20             = 4'h0;
assign OE_DATA_64_const_net_20             = 4'h0;
assign OE_DATA_65_const_net_20             = 4'h0;
assign OE_DATA_66_const_net_20             = 4'h0;
assign OE_DATA_67_const_net_20             = 4'h0;
assign OE_DATA_68_const_net_20             = 4'h0;
assign OE_DATA_69_const_net_20             = 4'h0;
assign OE_DATA_70_const_net_20             = 4'h0;
assign OE_DATA_71_const_net_20             = 4'h0;
assign OE_DATA_72_const_net_20             = 4'h0;
assign OE_DATA_73_const_net_20             = 4'h0;
assign OE_DATA_74_const_net_20             = 4'h0;
assign OE_DATA_75_const_net_20             = 4'h0;
assign OE_DATA_76_const_net_20             = 4'h0;
assign OE_DATA_77_const_net_20             = 4'h0;
assign OE_DATA_78_const_net_20             = 4'h0;
assign OE_DATA_79_const_net_20             = 4'h0;
assign OE_DATA_80_const_net_20             = 4'h0;
assign OE_DATA_81_const_net_20             = 4'h0;
assign OE_DATA_82_const_net_20             = 4'h0;
assign OE_DATA_83_const_net_20             = 4'h0;
assign OE_DATA_84_const_net_20             = 4'h0;
assign OE_DATA_85_const_net_20             = 4'h0;
assign OE_DATA_86_const_net_20             = 4'h0;
assign OE_DATA_87_const_net_20             = 4'h0;
assign OE_DATA_88_const_net_20             = 4'h0;
assign OE_DATA_89_const_net_20             = 4'h0;
assign OE_DATA_90_const_net_20             = 4'h0;
assign OE_DATA_91_const_net_20             = 4'h0;
assign OE_DATA_92_const_net_20             = 4'h0;
assign OE_DATA_93_const_net_20             = 4'h0;
assign OE_DATA_94_const_net_20             = 4'h0;
assign OE_DATA_95_const_net_20             = 4'h0;
assign OE_DATA_96_const_net_20             = 4'h0;
assign OE_DATA_97_const_net_20             = 4'h0;
assign OE_DATA_98_const_net_20             = 4'h0;
assign OE_DATA_99_const_net_20             = 4'h0;
assign OE_DATA_100_const_net_20            = 4'h0;
assign OE_DATA_101_const_net_20            = 4'h0;
assign OE_DATA_102_const_net_20            = 4'h0;
assign OE_DATA_103_const_net_20            = 4'h0;
assign OE_DATA_104_const_net_20            = 4'h0;
assign OE_DATA_105_const_net_20            = 4'h0;
assign OE_DATA_106_const_net_20            = 4'h0;
assign OE_DATA_107_const_net_20            = 4'h0;
assign OE_DATA_108_const_net_20            = 4'h0;
assign OE_DATA_109_const_net_20            = 4'h0;
assign OE_DATA_110_const_net_20            = 4'h0;
assign OE_DATA_111_const_net_20            = 4'h0;
assign OE_DATA_112_const_net_20            = 4'h0;
assign OE_DATA_113_const_net_20            = 4'h0;
assign OE_DATA_114_const_net_20            = 4'h0;
assign OE_DATA_115_const_net_20            = 4'h0;
assign OE_DATA_116_const_net_20            = 4'h0;
assign OE_DATA_117_const_net_20            = 4'h0;
assign OE_DATA_118_const_net_20            = 4'h0;
assign OE_DATA_119_const_net_20            = 4'h0;
assign OE_DATA_120_const_net_20            = 4'h0;
assign OE_DATA_121_const_net_20            = 4'h0;
assign OE_DATA_122_const_net_20            = 4'h0;
assign OE_DATA_123_const_net_20            = 4'h0;
assign OE_DATA_124_const_net_20            = 4'h0;
assign OE_DATA_125_const_net_20            = 4'h0;
assign OE_DATA_126_const_net_20            = 4'h0;
assign OE_DATA_127_const_net_20            = 4'h0;
assign TX_DATA_8_const_net_20              = 8'h00;
assign TX_DATA_9_const_net_20              = 8'h00;
assign TX_DATA_10_const_net_20             = 8'h00;
assign TX_DATA_11_const_net_20             = 8'h00;
assign TX_DATA_12_const_net_21             = 8'h00;
assign TX_DATA_13_const_net_21             = 8'h00;
assign TX_DATA_14_const_net_21             = 8'h00;
assign TX_DATA_15_const_net_21             = 8'h00;
assign TX_DATA_16_const_net_21             = 8'h00;
assign TX_DATA_17_const_net_21             = 8'h00;
assign TX_DATA_18_const_net_21             = 8'h00;
assign TX_DATA_19_const_net_21             = 8'h00;
assign TX_DATA_20_const_net_21             = 8'h00;
assign TX_DATA_21_const_net_21             = 8'h00;
assign TX_DATA_22_const_net_21             = 8'h00;
assign TX_DATA_23_const_net_21             = 8'h00;
assign TX_DATA_24_const_net_21             = 8'h00;
assign TX_DATA_25_const_net_21             = 8'h00;
assign TX_DATA_26_const_net_21             = 8'h00;
assign TX_DATA_27_const_net_21             = 8'h00;
assign TX_DATA_28_const_net_21             = 8'h00;
assign TX_DATA_29_const_net_21             = 8'h00;
assign TX_DATA_30_const_net_21             = 8'h00;
assign TX_DATA_31_const_net_21             = 8'h00;
assign TX_DATA_32_const_net_21             = 8'h00;
assign TX_DATA_33_const_net_21             = 8'h00;
assign TX_DATA_34_const_net_21             = 8'h00;
assign TX_DATA_35_const_net_21             = 8'h00;
assign TX_DATA_36_const_net_21             = 8'h00;
assign TX_DATA_37_const_net_21             = 8'h00;
assign TX_DATA_38_const_net_21             = 8'h00;
assign TX_DATA_39_const_net_21             = 8'h00;
assign TX_DATA_40_const_net_21             = 8'h00;
assign TX_DATA_41_const_net_21             = 8'h00;
assign TX_DATA_42_const_net_21             = 8'h00;
assign TX_DATA_43_const_net_21             = 8'h00;
assign TX_DATA_44_const_net_21             = 8'h00;
assign TX_DATA_45_const_net_21             = 8'h00;
assign TX_DATA_46_const_net_21             = 8'h00;
assign TX_DATA_47_const_net_21             = 8'h00;
assign TX_DATA_48_const_net_21             = 8'h00;
assign TX_DATA_49_const_net_21             = 8'h00;
assign TX_DATA_50_const_net_21             = 8'h00;
assign TX_DATA_51_const_net_21             = 8'h00;
assign TX_DATA_52_const_net_21             = 8'h00;
assign TX_DATA_53_const_net_21             = 8'h00;
assign TX_DATA_54_const_net_21             = 8'h00;
assign TX_DATA_55_const_net_21             = 8'h00;
assign TX_DATA_56_const_net_21             = 8'h00;
assign TX_DATA_57_const_net_21             = 8'h00;
assign TX_DATA_58_const_net_21             = 8'h00;
assign TX_DATA_59_const_net_21             = 8'h00;
assign TX_DATA_60_const_net_21             = 8'h00;
assign TX_DATA_61_const_net_21             = 8'h00;
assign TX_DATA_62_const_net_21             = 8'h00;
assign TX_DATA_63_const_net_21             = 8'h00;
assign TX_DATA_64_const_net_21             = 8'h00;
assign TX_DATA_65_const_net_21             = 8'h00;
assign TX_DATA_66_const_net_21             = 8'h00;
assign TX_DATA_67_const_net_21             = 8'h00;
assign TX_DATA_68_const_net_21             = 8'h00;
assign TX_DATA_69_const_net_21             = 8'h00;
assign TX_DATA_70_const_net_21             = 8'h00;
assign TX_DATA_71_const_net_21             = 8'h00;
assign TX_DATA_72_const_net_21             = 8'h00;
assign TX_DATA_73_const_net_21             = 8'h00;
assign TX_DATA_74_const_net_21             = 8'h00;
assign TX_DATA_75_const_net_21             = 8'h00;
assign TX_DATA_76_const_net_21             = 8'h00;
assign TX_DATA_77_const_net_21             = 8'h00;
assign TX_DATA_78_const_net_21             = 8'h00;
assign TX_DATA_79_const_net_21             = 8'h00;
assign TX_DATA_80_const_net_21             = 8'h00;
assign TX_DATA_81_const_net_21             = 8'h00;
assign TX_DATA_82_const_net_21             = 8'h00;
assign TX_DATA_83_const_net_21             = 8'h00;
assign TX_DATA_84_const_net_21             = 8'h00;
assign TX_DATA_85_const_net_21             = 8'h00;
assign TX_DATA_86_const_net_21             = 8'h00;
assign TX_DATA_87_const_net_21             = 8'h00;
assign TX_DATA_88_const_net_21             = 8'h00;
assign TX_DATA_89_const_net_21             = 8'h00;
assign TX_DATA_90_const_net_21             = 8'h00;
assign TX_DATA_91_const_net_21             = 8'h00;
assign TX_DATA_92_const_net_21             = 8'h00;
assign TX_DATA_93_const_net_21             = 8'h00;
assign TX_DATA_94_const_net_21             = 8'h00;
assign TX_DATA_95_const_net_21             = 8'h00;
assign TX_DATA_96_const_net_21             = 8'h00;
assign TX_DATA_97_const_net_21             = 8'h00;
assign TX_DATA_98_const_net_21             = 8'h00;
assign TX_DATA_99_const_net_21             = 8'h00;
assign TX_DATA_100_const_net_21            = 8'h00;
assign TX_DATA_101_const_net_21            = 8'h00;
assign TX_DATA_102_const_net_21            = 8'h00;
assign TX_DATA_103_const_net_21            = 8'h00;
assign TX_DATA_104_const_net_21            = 8'h00;
assign TX_DATA_105_const_net_21            = 8'h00;
assign TX_DATA_106_const_net_21            = 8'h00;
assign TX_DATA_107_const_net_21            = 8'h00;
assign TX_DATA_108_const_net_21            = 8'h00;
assign TX_DATA_109_const_net_21            = 8'h00;
assign TX_DATA_110_const_net_21            = 8'h00;
assign TX_DATA_111_const_net_21            = 8'h00;
assign TX_DATA_112_const_net_21            = 8'h00;
assign TX_DATA_113_const_net_21            = 8'h00;
assign TX_DATA_114_const_net_21            = 8'h00;
assign TX_DATA_115_const_net_21            = 8'h00;
assign TX_DATA_116_const_net_21            = 8'h00;
assign TX_DATA_117_const_net_21            = 8'h00;
assign TX_DATA_118_const_net_21            = 8'h00;
assign TX_DATA_119_const_net_21            = 8'h00;
assign TX_DATA_120_const_net_21            = 8'h00;
assign TX_DATA_121_const_net_21            = 8'h00;
assign TX_DATA_122_const_net_21            = 8'h00;
assign TX_DATA_123_const_net_21            = 8'h00;
assign TX_DATA_124_const_net_21            = 8'h00;
assign TX_DATA_125_const_net_21            = 8'h00;
assign TX_DATA_126_const_net_21            = 8'h00;
assign TX_DATA_127_const_net_21            = 8'h00;
assign OE_DATA_8_const_net_21              = 4'h0;
assign OE_DATA_9_const_net_21              = 4'h0;
assign OE_DATA_10_const_net_21             = 4'h0;
assign OE_DATA_11_const_net_21             = 4'h0;
assign OE_DATA_12_const_net_21             = 4'h0;
assign OE_DATA_13_const_net_21             = 4'h0;
assign OE_DATA_14_const_net_21             = 4'h0;
assign OE_DATA_15_const_net_21             = 4'h0;
assign OE_DATA_16_const_net_21             = 4'h0;
assign OE_DATA_17_const_net_21             = 4'h0;
assign OE_DATA_18_const_net_21             = 4'h0;
assign OE_DATA_19_const_net_21             = 4'h0;
assign OE_DATA_20_const_net_21             = 4'h0;
assign OE_DATA_21_const_net_21             = 4'h0;
assign OE_DATA_22_const_net_21             = 4'h0;
assign OE_DATA_23_const_net_21             = 4'h0;
assign OE_DATA_24_const_net_21             = 4'h0;
assign OE_DATA_25_const_net_21             = 4'h0;
assign OE_DATA_26_const_net_21             = 4'h0;
assign OE_DATA_27_const_net_21             = 4'h0;
assign OE_DATA_28_const_net_21             = 4'h0;
assign OE_DATA_29_const_net_21             = 4'h0;
assign OE_DATA_30_const_net_21             = 4'h0;
assign OE_DATA_31_const_net_21             = 4'h0;
assign OE_DATA_32_const_net_21             = 4'h0;
assign OE_DATA_33_const_net_21             = 4'h0;
assign OE_DATA_34_const_net_21             = 4'h0;
assign OE_DATA_35_const_net_21             = 4'h0;
assign OE_DATA_36_const_net_21             = 4'h0;
assign OE_DATA_37_const_net_21             = 4'h0;
assign OE_DATA_38_const_net_21             = 4'h0;
assign OE_DATA_39_const_net_21             = 4'h0;
assign OE_DATA_40_const_net_21             = 4'h0;
assign OE_DATA_41_const_net_21             = 4'h0;
assign OE_DATA_42_const_net_21             = 4'h0;
assign OE_DATA_43_const_net_21             = 4'h0;
assign OE_DATA_44_const_net_21             = 4'h0;
assign OE_DATA_45_const_net_21             = 4'h0;
assign OE_DATA_46_const_net_21             = 4'h0;
assign OE_DATA_47_const_net_21             = 4'h0;
assign OE_DATA_48_const_net_21             = 4'h0;
assign OE_DATA_49_const_net_21             = 4'h0;
assign OE_DATA_50_const_net_21             = 4'h0;
assign OE_DATA_51_const_net_21             = 4'h0;
assign OE_DATA_52_const_net_21             = 4'h0;
assign OE_DATA_53_const_net_21             = 4'h0;
assign OE_DATA_54_const_net_21             = 4'h0;
assign OE_DATA_55_const_net_21             = 4'h0;
assign OE_DATA_56_const_net_21             = 4'h0;
assign OE_DATA_57_const_net_21             = 4'h0;
assign OE_DATA_58_const_net_21             = 4'h0;
assign OE_DATA_59_const_net_21             = 4'h0;
assign OE_DATA_60_const_net_21             = 4'h0;
assign OE_DATA_61_const_net_21             = 4'h0;
assign OE_DATA_62_const_net_21             = 4'h0;
assign OE_DATA_63_const_net_21             = 4'h0;
assign OE_DATA_64_const_net_21             = 4'h0;
assign OE_DATA_65_const_net_21             = 4'h0;
assign OE_DATA_66_const_net_21             = 4'h0;
assign OE_DATA_67_const_net_21             = 4'h0;
assign OE_DATA_68_const_net_21             = 4'h0;
assign OE_DATA_69_const_net_21             = 4'h0;
assign OE_DATA_70_const_net_21             = 4'h0;
assign OE_DATA_71_const_net_21             = 4'h0;
assign OE_DATA_72_const_net_21             = 4'h0;
assign OE_DATA_73_const_net_21             = 4'h0;
assign OE_DATA_74_const_net_21             = 4'h0;
assign OE_DATA_75_const_net_21             = 4'h0;
assign OE_DATA_76_const_net_21             = 4'h0;
assign OE_DATA_77_const_net_21             = 4'h0;
assign OE_DATA_78_const_net_21             = 4'h0;
assign OE_DATA_79_const_net_21             = 4'h0;
assign OE_DATA_80_const_net_21             = 4'h0;
assign OE_DATA_81_const_net_21             = 4'h0;
assign OE_DATA_82_const_net_21             = 4'h0;
assign OE_DATA_83_const_net_21             = 4'h0;
assign OE_DATA_84_const_net_21             = 4'h0;
assign OE_DATA_85_const_net_21             = 4'h0;
assign OE_DATA_86_const_net_21             = 4'h0;
assign OE_DATA_87_const_net_21             = 4'h0;
assign OE_DATA_88_const_net_21             = 4'h0;
assign OE_DATA_89_const_net_21             = 4'h0;
assign OE_DATA_90_const_net_21             = 4'h0;
assign OE_DATA_91_const_net_21             = 4'h0;
assign OE_DATA_92_const_net_21             = 4'h0;
assign OE_DATA_93_const_net_21             = 4'h0;
assign OE_DATA_94_const_net_21             = 4'h0;
assign OE_DATA_95_const_net_21             = 4'h0;
assign OE_DATA_96_const_net_21             = 4'h0;
assign OE_DATA_97_const_net_21             = 4'h0;
assign OE_DATA_98_const_net_21             = 4'h0;
assign OE_DATA_99_const_net_21             = 4'h0;
assign OE_DATA_100_const_net_21            = 4'h0;
assign OE_DATA_101_const_net_21            = 4'h0;
assign OE_DATA_102_const_net_21            = 4'h0;
assign OE_DATA_103_const_net_21            = 4'h0;
assign OE_DATA_104_const_net_21            = 4'h0;
assign OE_DATA_105_const_net_21            = 4'h0;
assign OE_DATA_106_const_net_21            = 4'h0;
assign OE_DATA_107_const_net_21            = 4'h0;
assign OE_DATA_108_const_net_21            = 4'h0;
assign OE_DATA_109_const_net_21            = 4'h0;
assign OE_DATA_110_const_net_21            = 4'h0;
assign OE_DATA_111_const_net_21            = 4'h0;
assign OE_DATA_112_const_net_21            = 4'h0;
assign OE_DATA_113_const_net_21            = 4'h0;
assign OE_DATA_114_const_net_21            = 4'h0;
assign OE_DATA_115_const_net_21            = 4'h0;
assign OE_DATA_116_const_net_21            = 4'h0;
assign OE_DATA_117_const_net_21            = 4'h0;
assign OE_DATA_118_const_net_21            = 4'h0;
assign OE_DATA_119_const_net_21            = 4'h0;
assign OE_DATA_120_const_net_21            = 4'h0;
assign OE_DATA_121_const_net_21            = 4'h0;
assign OE_DATA_122_const_net_21            = 4'h0;
assign OE_DATA_123_const_net_21            = 4'h0;
assign OE_DATA_124_const_net_21            = 4'h0;
assign OE_DATA_125_const_net_21            = 4'h0;
assign OE_DATA_126_const_net_21            = 4'h0;
assign OE_DATA_127_const_net_21            = 4'h0;
assign PAD_I_const_net_4                   = 8'h00;
assign PAD_N_const_net_4                   = 8'h00;
assign PAD_I_N_const_net_4                 = 8'h00;
assign TX_DATA_1_const_net_17              = 8'h00;
assign TX_DATA_2_const_net_19              = 8'h00;
assign TX_DATA_3_const_net_19              = 8'h00;
assign TX_DATA_4_const_net_19              = 8'h00;
assign TX_DATA_5_const_net_19              = 8'h00;
assign TX_DATA_6_const_net_19              = 8'h00;
assign TX_DATA_7_const_net_19              = 8'h00;
assign TX_DATA_8_const_net_21              = 8'h00;
assign TX_DATA_9_const_net_21              = 8'h00;
assign TX_DATA_10_const_net_21             = 8'h00;
assign TX_DATA_11_const_net_21             = 8'h00;
assign TX_DATA_12_const_net_22             = 8'h00;
assign TX_DATA_13_const_net_22             = 8'h00;
assign TX_DATA_14_const_net_22             = 8'h00;
assign TX_DATA_15_const_net_22             = 8'h00;
assign TX_DATA_16_const_net_22             = 8'h00;
assign TX_DATA_17_const_net_22             = 8'h00;
assign TX_DATA_18_const_net_22             = 8'h00;
assign TX_DATA_19_const_net_22             = 8'h00;
assign TX_DATA_20_const_net_22             = 8'h00;
assign TX_DATA_21_const_net_22             = 8'h00;
assign TX_DATA_22_const_net_22             = 8'h00;
assign TX_DATA_23_const_net_22             = 8'h00;
assign TX_DATA_24_const_net_22             = 8'h00;
assign TX_DATA_25_const_net_22             = 8'h00;
assign TX_DATA_26_const_net_22             = 8'h00;
assign TX_DATA_27_const_net_22             = 8'h00;
assign TX_DATA_28_const_net_22             = 8'h00;
assign TX_DATA_29_const_net_22             = 8'h00;
assign TX_DATA_30_const_net_22             = 8'h00;
assign TX_DATA_31_const_net_22             = 8'h00;
assign TX_DATA_32_const_net_22             = 8'h00;
assign TX_DATA_33_const_net_22             = 8'h00;
assign TX_DATA_34_const_net_22             = 8'h00;
assign TX_DATA_35_const_net_22             = 8'h00;
assign TX_DATA_36_const_net_22             = 8'h00;
assign TX_DATA_37_const_net_22             = 8'h00;
assign TX_DATA_38_const_net_22             = 8'h00;
assign TX_DATA_39_const_net_22             = 8'h00;
assign TX_DATA_40_const_net_22             = 8'h00;
assign TX_DATA_41_const_net_22             = 8'h00;
assign TX_DATA_42_const_net_22             = 8'h00;
assign TX_DATA_43_const_net_22             = 8'h00;
assign TX_DATA_44_const_net_22             = 8'h00;
assign TX_DATA_45_const_net_22             = 8'h00;
assign TX_DATA_46_const_net_22             = 8'h00;
assign TX_DATA_47_const_net_22             = 8'h00;
assign TX_DATA_48_const_net_22             = 8'h00;
assign TX_DATA_49_const_net_22             = 8'h00;
assign TX_DATA_50_const_net_22             = 8'h00;
assign TX_DATA_51_const_net_22             = 8'h00;
assign TX_DATA_52_const_net_22             = 8'h00;
assign TX_DATA_53_const_net_22             = 8'h00;
assign TX_DATA_54_const_net_22             = 8'h00;
assign TX_DATA_55_const_net_22             = 8'h00;
assign TX_DATA_56_const_net_22             = 8'h00;
assign TX_DATA_57_const_net_22             = 8'h00;
assign TX_DATA_58_const_net_22             = 8'h00;
assign TX_DATA_59_const_net_22             = 8'h00;
assign TX_DATA_60_const_net_22             = 8'h00;
assign TX_DATA_61_const_net_22             = 8'h00;
assign TX_DATA_62_const_net_22             = 8'h00;
assign TX_DATA_63_const_net_22             = 8'h00;
assign TX_DATA_64_const_net_22             = 8'h00;
assign TX_DATA_65_const_net_22             = 8'h00;
assign TX_DATA_66_const_net_22             = 8'h00;
assign TX_DATA_67_const_net_22             = 8'h00;
assign TX_DATA_68_const_net_22             = 8'h00;
assign TX_DATA_69_const_net_22             = 8'h00;
assign TX_DATA_70_const_net_22             = 8'h00;
assign TX_DATA_71_const_net_22             = 8'h00;
assign TX_DATA_72_const_net_22             = 8'h00;
assign TX_DATA_73_const_net_22             = 8'h00;
assign TX_DATA_74_const_net_22             = 8'h00;
assign TX_DATA_75_const_net_22             = 8'h00;
assign TX_DATA_76_const_net_22             = 8'h00;
assign TX_DATA_77_const_net_22             = 8'h00;
assign TX_DATA_78_const_net_22             = 8'h00;
assign TX_DATA_79_const_net_22             = 8'h00;
assign TX_DATA_80_const_net_22             = 8'h00;
assign TX_DATA_81_const_net_22             = 8'h00;
assign TX_DATA_82_const_net_22             = 8'h00;
assign TX_DATA_83_const_net_22             = 8'h00;
assign TX_DATA_84_const_net_22             = 8'h00;
assign TX_DATA_85_const_net_22             = 8'h00;
assign TX_DATA_86_const_net_22             = 8'h00;
assign TX_DATA_87_const_net_22             = 8'h00;
assign TX_DATA_88_const_net_22             = 8'h00;
assign TX_DATA_89_const_net_22             = 8'h00;
assign TX_DATA_90_const_net_22             = 8'h00;
assign TX_DATA_91_const_net_22             = 8'h00;
assign TX_DATA_92_const_net_22             = 8'h00;
assign TX_DATA_93_const_net_22             = 8'h00;
assign TX_DATA_94_const_net_22             = 8'h00;
assign TX_DATA_95_const_net_22             = 8'h00;
assign TX_DATA_96_const_net_22             = 8'h00;
assign TX_DATA_97_const_net_22             = 8'h00;
assign TX_DATA_98_const_net_22             = 8'h00;
assign TX_DATA_99_const_net_22             = 8'h00;
assign TX_DATA_100_const_net_22            = 8'h00;
assign TX_DATA_101_const_net_22            = 8'h00;
assign TX_DATA_102_const_net_22            = 8'h00;
assign TX_DATA_103_const_net_22            = 8'h00;
assign TX_DATA_104_const_net_22            = 8'h00;
assign TX_DATA_105_const_net_22            = 8'h00;
assign TX_DATA_106_const_net_22            = 8'h00;
assign TX_DATA_107_const_net_22            = 8'h00;
assign TX_DATA_108_const_net_22            = 8'h00;
assign TX_DATA_109_const_net_22            = 8'h00;
assign TX_DATA_110_const_net_22            = 8'h00;
assign TX_DATA_111_const_net_22            = 8'h00;
assign TX_DATA_112_const_net_22            = 8'h00;
assign TX_DATA_113_const_net_22            = 8'h00;
assign TX_DATA_114_const_net_22            = 8'h00;
assign TX_DATA_115_const_net_22            = 8'h00;
assign TX_DATA_116_const_net_22            = 8'h00;
assign TX_DATA_117_const_net_22            = 8'h00;
assign TX_DATA_118_const_net_22            = 8'h00;
assign TX_DATA_119_const_net_22            = 8'h00;
assign TX_DATA_120_const_net_22            = 8'h00;
assign TX_DATA_121_const_net_22            = 8'h00;
assign TX_DATA_122_const_net_22            = 8'h00;
assign TX_DATA_123_const_net_22            = 8'h00;
assign TX_DATA_124_const_net_22            = 8'h00;
assign TX_DATA_125_const_net_22            = 8'h00;
assign TX_DATA_126_const_net_22            = 8'h00;
assign TX_DATA_127_const_net_22            = 8'h00;
assign OE_DATA_1_const_net_20              = 4'h0;
assign OE_DATA_2_const_net_20              = 4'h0;
assign OE_DATA_3_const_net_20              = 4'h0;
assign OE_DATA_4_const_net_20              = 4'h0;
assign OE_DATA_5_const_net_20              = 4'h0;
assign OE_DATA_6_const_net_20              = 4'h0;
assign OE_DATA_7_const_net_20              = 4'h0;
assign OE_DATA_8_const_net_22              = 4'h0;
assign OE_DATA_9_const_net_22              = 4'h0;
assign OE_DATA_10_const_net_22             = 4'h0;
assign OE_DATA_11_const_net_22             = 4'h0;
assign OE_DATA_12_const_net_22             = 4'h0;
assign OE_DATA_13_const_net_22             = 4'h0;
assign OE_DATA_14_const_net_22             = 4'h0;
assign OE_DATA_15_const_net_22             = 4'h0;
assign OE_DATA_16_const_net_22             = 4'h0;
assign OE_DATA_17_const_net_22             = 4'h0;
assign OE_DATA_18_const_net_22             = 4'h0;
assign OE_DATA_19_const_net_22             = 4'h0;
assign OE_DATA_20_const_net_22             = 4'h0;
assign OE_DATA_21_const_net_22             = 4'h0;
assign OE_DATA_22_const_net_22             = 4'h0;
assign OE_DATA_23_const_net_22             = 4'h0;
assign OE_DATA_24_const_net_22             = 4'h0;
assign OE_DATA_25_const_net_22             = 4'h0;
assign OE_DATA_26_const_net_22             = 4'h0;
assign OE_DATA_27_const_net_22             = 4'h0;
assign OE_DATA_28_const_net_22             = 4'h0;
assign OE_DATA_29_const_net_22             = 4'h0;
assign OE_DATA_30_const_net_22             = 4'h0;
assign OE_DATA_31_const_net_22             = 4'h0;
assign OE_DATA_32_const_net_22             = 4'h0;
assign OE_DATA_33_const_net_22             = 4'h0;
assign OE_DATA_34_const_net_22             = 4'h0;
assign OE_DATA_35_const_net_22             = 4'h0;
assign OE_DATA_36_const_net_22             = 4'h0;
assign OE_DATA_37_const_net_22             = 4'h0;
assign OE_DATA_38_const_net_22             = 4'h0;
assign OE_DATA_39_const_net_22             = 4'h0;
assign OE_DATA_40_const_net_22             = 4'h0;
assign OE_DATA_41_const_net_22             = 4'h0;
assign OE_DATA_42_const_net_22             = 4'h0;
assign OE_DATA_43_const_net_22             = 4'h0;
assign OE_DATA_44_const_net_22             = 4'h0;
assign OE_DATA_45_const_net_22             = 4'h0;
assign OE_DATA_46_const_net_22             = 4'h0;
assign OE_DATA_47_const_net_22             = 4'h0;
assign OE_DATA_48_const_net_22             = 4'h0;
assign OE_DATA_49_const_net_22             = 4'h0;
assign OE_DATA_50_const_net_22             = 4'h0;
assign OE_DATA_51_const_net_22             = 4'h0;
assign OE_DATA_52_const_net_22             = 4'h0;
assign OE_DATA_53_const_net_22             = 4'h0;
assign OE_DATA_54_const_net_22             = 4'h0;
assign OE_DATA_55_const_net_22             = 4'h0;
assign OE_DATA_56_const_net_22             = 4'h0;
assign OE_DATA_57_const_net_22             = 4'h0;
assign OE_DATA_58_const_net_22             = 4'h0;
assign OE_DATA_59_const_net_22             = 4'h0;
assign OE_DATA_60_const_net_22             = 4'h0;
assign OE_DATA_61_const_net_22             = 4'h0;
assign OE_DATA_62_const_net_22             = 4'h0;
assign OE_DATA_63_const_net_22             = 4'h0;
assign OE_DATA_64_const_net_22             = 4'h0;
assign OE_DATA_65_const_net_22             = 4'h0;
assign OE_DATA_66_const_net_22             = 4'h0;
assign OE_DATA_67_const_net_22             = 4'h0;
assign OE_DATA_68_const_net_22             = 4'h0;
assign OE_DATA_69_const_net_22             = 4'h0;
assign OE_DATA_70_const_net_22             = 4'h0;
assign OE_DATA_71_const_net_22             = 4'h0;
assign OE_DATA_72_const_net_22             = 4'h0;
assign OE_DATA_73_const_net_22             = 4'h0;
assign OE_DATA_74_const_net_22             = 4'h0;
assign OE_DATA_75_const_net_22             = 4'h0;
assign OE_DATA_76_const_net_22             = 4'h0;
assign OE_DATA_77_const_net_22             = 4'h0;
assign OE_DATA_78_const_net_22             = 4'h0;
assign OE_DATA_79_const_net_22             = 4'h0;
assign OE_DATA_80_const_net_22             = 4'h0;
assign OE_DATA_81_const_net_22             = 4'h0;
assign OE_DATA_82_const_net_22             = 4'h0;
assign OE_DATA_83_const_net_22             = 4'h0;
assign OE_DATA_84_const_net_22             = 4'h0;
assign OE_DATA_85_const_net_22             = 4'h0;
assign OE_DATA_86_const_net_22             = 4'h0;
assign OE_DATA_87_const_net_22             = 4'h0;
assign OE_DATA_88_const_net_22             = 4'h0;
assign OE_DATA_89_const_net_22             = 4'h0;
assign OE_DATA_90_const_net_22             = 4'h0;
assign OE_DATA_91_const_net_22             = 4'h0;
assign OE_DATA_92_const_net_22             = 4'h0;
assign OE_DATA_93_const_net_22             = 4'h0;
assign OE_DATA_94_const_net_22             = 4'h0;
assign OE_DATA_95_const_net_22             = 4'h0;
assign OE_DATA_96_const_net_22             = 4'h0;
assign OE_DATA_97_const_net_22             = 4'h0;
assign OE_DATA_98_const_net_22             = 4'h0;
assign OE_DATA_99_const_net_22             = 4'h0;
assign OE_DATA_100_const_net_22            = 4'h0;
assign OE_DATA_101_const_net_22            = 4'h0;
assign OE_DATA_102_const_net_22            = 4'h0;
assign OE_DATA_103_const_net_22            = 4'h0;
assign OE_DATA_104_const_net_22            = 4'h0;
assign OE_DATA_105_const_net_22            = 4'h0;
assign OE_DATA_106_const_net_22            = 4'h0;
assign OE_DATA_107_const_net_22            = 4'h0;
assign OE_DATA_108_const_net_22            = 4'h0;
assign OE_DATA_109_const_net_22            = 4'h0;
assign OE_DATA_110_const_net_22            = 4'h0;
assign OE_DATA_111_const_net_22            = 4'h0;
assign OE_DATA_112_const_net_22            = 4'h0;
assign OE_DATA_113_const_net_22            = 4'h0;
assign OE_DATA_114_const_net_22            = 4'h0;
assign OE_DATA_115_const_net_22            = 4'h0;
assign OE_DATA_116_const_net_22            = 4'h0;
assign OE_DATA_117_const_net_22            = 4'h0;
assign OE_DATA_118_const_net_22            = 4'h0;
assign OE_DATA_119_const_net_22            = 4'h0;
assign OE_DATA_120_const_net_22            = 4'h0;
assign OE_DATA_121_const_net_22            = 4'h0;
assign OE_DATA_122_const_net_22            = 4'h0;
assign OE_DATA_123_const_net_22            = 4'h0;
assign OE_DATA_124_const_net_22            = 4'h0;
assign OE_DATA_125_const_net_22            = 4'h0;
assign OE_DATA_126_const_net_22            = 4'h0;
assign OE_DATA_127_const_net_22            = 4'h0;
assign RX_DQS_90_const_net_17              = 2'h0;
assign FIFO_WR_PTR_const_net_18            = 3'h0;
assign FIFO_RD_PTR_const_net_18            = 3'h0;
assign EYE_MONITOR_LANE_WIDTH_const_net_19 = 3'h0;
assign TX_DATA_1_const_net_18              = 2'h0;
assign TX_DATA_2_const_net_20              = 2'h0;
assign TX_DATA_3_const_net_20              = 2'h0;
assign TX_DATA_4_const_net_20              = 2'h0;
assign TX_DATA_5_const_net_20              = 2'h0;
assign TX_DATA_6_const_net_20              = 2'h0;
assign TX_DATA_7_const_net_20              = 2'h0;
assign TX_DATA_8_const_net_22              = 2'h0;
assign TX_DATA_9_const_net_22              = 2'h0;
assign TX_DATA_10_const_net_22             = 2'h0;
assign TX_DATA_11_const_net_22             = 2'h0;
assign TX_DATA_12_const_net_23             = 2'h0;
assign TX_DATA_13_const_net_23             = 2'h0;
assign TX_DATA_14_const_net_23             = 2'h0;
assign TX_DATA_15_const_net_23             = 2'h0;
assign TX_DATA_16_const_net_23             = 2'h0;
assign TX_DATA_17_const_net_23             = 2'h0;
assign TX_DATA_18_const_net_23             = 2'h0;
assign TX_DATA_19_const_net_23             = 2'h0;
assign TX_DATA_20_const_net_23             = 2'h0;
assign TX_DATA_21_const_net_23             = 2'h0;
assign TX_DATA_22_const_net_23             = 2'h0;
assign TX_DATA_23_const_net_23             = 2'h0;
assign TX_DATA_24_const_net_23             = 2'h0;
assign TX_DATA_25_const_net_23             = 2'h0;
assign TX_DATA_26_const_net_23             = 2'h0;
assign TX_DATA_27_const_net_23             = 2'h0;
assign TX_DATA_28_const_net_23             = 2'h0;
assign TX_DATA_29_const_net_23             = 2'h0;
assign TX_DATA_30_const_net_23             = 2'h0;
assign TX_DATA_31_const_net_23             = 2'h0;
assign TX_DATA_32_const_net_23             = 2'h0;
assign TX_DATA_33_const_net_23             = 2'h0;
assign TX_DATA_34_const_net_23             = 2'h0;
assign TX_DATA_35_const_net_23             = 2'h0;
assign TX_DATA_36_const_net_23             = 2'h0;
assign TX_DATA_37_const_net_23             = 2'h0;
assign TX_DATA_38_const_net_23             = 2'h0;
assign TX_DATA_39_const_net_23             = 2'h0;
assign TX_DATA_40_const_net_23             = 2'h0;
assign TX_DATA_41_const_net_23             = 2'h0;
assign TX_DATA_42_const_net_23             = 2'h0;
assign TX_DATA_43_const_net_23             = 2'h0;
assign TX_DATA_44_const_net_23             = 2'h0;
assign TX_DATA_45_const_net_23             = 2'h0;
assign TX_DATA_46_const_net_23             = 2'h0;
assign TX_DATA_47_const_net_23             = 2'h0;
assign TX_DATA_48_const_net_23             = 2'h0;
assign TX_DATA_49_const_net_23             = 2'h0;
assign TX_DATA_50_const_net_23             = 2'h0;
assign TX_DATA_51_const_net_23             = 2'h0;
assign TX_DATA_52_const_net_23             = 2'h0;
assign TX_DATA_53_const_net_23             = 2'h0;
assign TX_DATA_54_const_net_23             = 2'h0;
assign TX_DATA_55_const_net_23             = 2'h0;
assign TX_DATA_56_const_net_23             = 2'h0;
assign TX_DATA_57_const_net_23             = 2'h0;
assign TX_DATA_58_const_net_23             = 2'h0;
assign TX_DATA_59_const_net_23             = 2'h0;
assign TX_DATA_60_const_net_23             = 2'h0;
assign TX_DATA_61_const_net_23             = 2'h0;
assign TX_DATA_62_const_net_23             = 2'h0;
assign TX_DATA_63_const_net_23             = 2'h0;
assign TX_DATA_64_const_net_23             = 2'h0;
assign TX_DATA_65_const_net_23             = 2'h0;
assign TX_DATA_66_const_net_23             = 2'h0;
assign TX_DATA_67_const_net_23             = 2'h0;
assign TX_DATA_68_const_net_23             = 2'h0;
assign TX_DATA_69_const_net_23             = 2'h0;
assign TX_DATA_70_const_net_23             = 2'h0;
assign TX_DATA_71_const_net_23             = 2'h0;
assign TX_DATA_72_const_net_23             = 2'h0;
assign TX_DATA_73_const_net_23             = 2'h0;
assign TX_DATA_74_const_net_23             = 2'h0;
assign TX_DATA_75_const_net_23             = 2'h0;
assign TX_DATA_76_const_net_23             = 2'h0;
assign TX_DATA_77_const_net_23             = 2'h0;
assign TX_DATA_78_const_net_23             = 2'h0;
assign TX_DATA_79_const_net_23             = 2'h0;
assign TX_DATA_80_const_net_23             = 2'h0;
assign TX_DATA_81_const_net_23             = 2'h0;
assign TX_DATA_82_const_net_23             = 2'h0;
assign TX_DATA_83_const_net_23             = 2'h0;
assign TX_DATA_84_const_net_23             = 2'h0;
assign TX_DATA_85_const_net_23             = 2'h0;
assign TX_DATA_86_const_net_23             = 2'h0;
assign TX_DATA_87_const_net_23             = 2'h0;
assign TX_DATA_88_const_net_23             = 2'h0;
assign TX_DATA_89_const_net_23             = 2'h0;
assign TX_DATA_90_const_net_23             = 2'h0;
assign TX_DATA_91_const_net_23             = 2'h0;
assign TX_DATA_92_const_net_23             = 2'h0;
assign TX_DATA_93_const_net_23             = 2'h0;
assign TX_DATA_94_const_net_23             = 2'h0;
assign TX_DATA_95_const_net_23             = 2'h0;
assign TX_DATA_96_const_net_23             = 2'h0;
assign TX_DATA_97_const_net_23             = 2'h0;
assign TX_DATA_98_const_net_23             = 2'h0;
assign TX_DATA_99_const_net_23             = 2'h0;
assign TX_DATA_100_const_net_23            = 2'h0;
assign TX_DATA_101_const_net_23            = 2'h0;
assign TX_DATA_102_const_net_23            = 2'h0;
assign TX_DATA_103_const_net_23            = 2'h0;
assign TX_DATA_104_const_net_23            = 2'h0;
assign TX_DATA_105_const_net_23            = 2'h0;
assign TX_DATA_106_const_net_23            = 2'h0;
assign TX_DATA_107_const_net_23            = 2'h0;
assign TX_DATA_108_const_net_23            = 2'h0;
assign TX_DATA_109_const_net_23            = 2'h0;
assign TX_DATA_110_const_net_23            = 2'h0;
assign TX_DATA_111_const_net_23            = 2'h0;
assign TX_DATA_112_const_net_23            = 2'h0;
assign TX_DATA_113_const_net_23            = 2'h0;
assign TX_DATA_114_const_net_23            = 2'h0;
assign TX_DATA_115_const_net_23            = 2'h0;
assign TX_DATA_116_const_net_23            = 2'h0;
assign TX_DATA_117_const_net_23            = 2'h0;
assign TX_DATA_118_const_net_23            = 2'h0;
assign TX_DATA_119_const_net_23            = 2'h0;
assign TX_DATA_120_const_net_23            = 2'h0;
assign TX_DATA_121_const_net_23            = 2'h0;
assign TX_DATA_122_const_net_23            = 2'h0;
assign TX_DATA_123_const_net_23            = 2'h0;
assign TX_DATA_124_const_net_23            = 2'h0;
assign TX_DATA_125_const_net_23            = 2'h0;
assign TX_DATA_126_const_net_23            = 2'h0;
assign TX_DATA_127_const_net_23            = 2'h0;
assign OE_DATA_1_const_net_21              = 2'h0;
assign OE_DATA_2_const_net_21              = 2'h0;
assign OE_DATA_3_const_net_21              = 2'h0;
assign OE_DATA_4_const_net_21              = 2'h0;
assign OE_DATA_5_const_net_21              = 2'h0;
assign OE_DATA_6_const_net_21              = 2'h0;
assign OE_DATA_7_const_net_21              = 2'h0;
assign OE_DATA_8_const_net_23              = 2'h0;
assign OE_DATA_9_const_net_23              = 2'h0;
assign OE_DATA_10_const_net_23             = 2'h0;
assign OE_DATA_11_const_net_23             = 2'h0;
assign OE_DATA_12_const_net_23             = 2'h0;
assign OE_DATA_13_const_net_23             = 2'h0;
assign OE_DATA_14_const_net_23             = 2'h0;
assign OE_DATA_15_const_net_23             = 2'h0;
assign OE_DATA_16_const_net_23             = 2'h0;
assign OE_DATA_17_const_net_23             = 2'h0;
assign OE_DATA_18_const_net_23             = 2'h0;
assign OE_DATA_19_const_net_23             = 2'h0;
assign OE_DATA_20_const_net_23             = 2'h0;
assign OE_DATA_21_const_net_23             = 2'h0;
assign OE_DATA_22_const_net_23             = 2'h0;
assign OE_DATA_23_const_net_23             = 2'h0;
assign OE_DATA_24_const_net_23             = 2'h0;
assign OE_DATA_25_const_net_23             = 2'h0;
assign OE_DATA_26_const_net_23             = 2'h0;
assign OE_DATA_27_const_net_23             = 2'h0;
assign OE_DATA_28_const_net_23             = 2'h0;
assign OE_DATA_29_const_net_23             = 2'h0;
assign OE_DATA_30_const_net_23             = 2'h0;
assign OE_DATA_31_const_net_23             = 2'h0;
assign OE_DATA_32_const_net_23             = 2'h0;
assign OE_DATA_33_const_net_23             = 2'h0;
assign OE_DATA_34_const_net_23             = 2'h0;
assign OE_DATA_35_const_net_23             = 2'h0;
assign OE_DATA_36_const_net_23             = 2'h0;
assign OE_DATA_37_const_net_23             = 2'h0;
assign OE_DATA_38_const_net_23             = 2'h0;
assign OE_DATA_39_const_net_23             = 2'h0;
assign OE_DATA_40_const_net_23             = 2'h0;
assign OE_DATA_41_const_net_23             = 2'h0;
assign OE_DATA_42_const_net_23             = 2'h0;
assign OE_DATA_43_const_net_23             = 2'h0;
assign OE_DATA_44_const_net_23             = 2'h0;
assign OE_DATA_45_const_net_23             = 2'h0;
assign OE_DATA_46_const_net_23             = 2'h0;
assign OE_DATA_47_const_net_23             = 2'h0;
assign OE_DATA_48_const_net_23             = 2'h0;
assign OE_DATA_49_const_net_23             = 2'h0;
assign OE_DATA_50_const_net_23             = 2'h0;
assign OE_DATA_51_const_net_23             = 2'h0;
assign OE_DATA_52_const_net_23             = 2'h0;
assign OE_DATA_53_const_net_23             = 2'h0;
assign OE_DATA_54_const_net_23             = 2'h0;
assign OE_DATA_55_const_net_23             = 2'h0;
assign OE_DATA_56_const_net_23             = 2'h0;
assign OE_DATA_57_const_net_23             = 2'h0;
assign OE_DATA_58_const_net_23             = 2'h0;
assign OE_DATA_59_const_net_23             = 2'h0;
assign OE_DATA_60_const_net_23             = 2'h0;
assign OE_DATA_61_const_net_23             = 2'h0;
assign OE_DATA_62_const_net_23             = 2'h0;
assign OE_DATA_63_const_net_23             = 2'h0;
assign OE_DATA_64_const_net_23             = 2'h0;
assign OE_DATA_65_const_net_23             = 2'h0;
assign OE_DATA_66_const_net_23             = 2'h0;
assign OE_DATA_67_const_net_23             = 2'h0;
assign OE_DATA_68_const_net_23             = 2'h0;
assign OE_DATA_69_const_net_23             = 2'h0;
assign OE_DATA_70_const_net_23             = 2'h0;
assign OE_DATA_71_const_net_23             = 2'h0;
assign OE_DATA_72_const_net_23             = 2'h0;
assign OE_DATA_73_const_net_23             = 2'h0;
assign OE_DATA_74_const_net_23             = 2'h0;
assign OE_DATA_75_const_net_23             = 2'h0;
assign OE_DATA_76_const_net_23             = 2'h0;
assign OE_DATA_77_const_net_23             = 2'h0;
assign OE_DATA_78_const_net_23             = 2'h0;
assign OE_DATA_79_const_net_23             = 2'h0;
assign OE_DATA_80_const_net_23             = 2'h0;
assign OE_DATA_81_const_net_23             = 2'h0;
assign OE_DATA_82_const_net_23             = 2'h0;
assign OE_DATA_83_const_net_23             = 2'h0;
assign OE_DATA_84_const_net_23             = 2'h0;
assign OE_DATA_85_const_net_23             = 2'h0;
assign OE_DATA_86_const_net_23             = 2'h0;
assign OE_DATA_87_const_net_23             = 2'h0;
assign OE_DATA_88_const_net_23             = 2'h0;
assign OE_DATA_89_const_net_23             = 2'h0;
assign OE_DATA_90_const_net_23             = 2'h0;
assign OE_DATA_91_const_net_23             = 2'h0;
assign OE_DATA_92_const_net_23             = 2'h0;
assign OE_DATA_93_const_net_23             = 2'h0;
assign OE_DATA_94_const_net_23             = 2'h0;
assign OE_DATA_95_const_net_23             = 2'h0;
assign OE_DATA_96_const_net_23             = 2'h0;
assign OE_DATA_97_const_net_23             = 2'h0;
assign OE_DATA_98_const_net_23             = 2'h0;
assign OE_DATA_99_const_net_23             = 2'h0;
assign OE_DATA_100_const_net_23            = 2'h0;
assign OE_DATA_101_const_net_23            = 2'h0;
assign OE_DATA_102_const_net_23            = 2'h0;
assign OE_DATA_103_const_net_23            = 2'h0;
assign OE_DATA_104_const_net_23            = 2'h0;
assign OE_DATA_105_const_net_23            = 2'h0;
assign OE_DATA_106_const_net_23            = 2'h0;
assign OE_DATA_107_const_net_23            = 2'h0;
assign OE_DATA_108_const_net_23            = 2'h0;
assign OE_DATA_109_const_net_23            = 2'h0;
assign OE_DATA_110_const_net_23            = 2'h0;
assign OE_DATA_111_const_net_23            = 2'h0;
assign OE_DATA_112_const_net_23            = 2'h0;
assign OE_DATA_113_const_net_23            = 2'h0;
assign OE_DATA_114_const_net_23            = 2'h0;
assign OE_DATA_115_const_net_23            = 2'h0;
assign OE_DATA_116_const_net_23            = 2'h0;
assign OE_DATA_117_const_net_23            = 2'h0;
assign OE_DATA_118_const_net_23            = 2'h0;
assign OE_DATA_119_const_net_23            = 2'h0;
assign OE_DATA_120_const_net_23            = 2'h0;
assign OE_DATA_121_const_net_23            = 2'h0;
assign OE_DATA_122_const_net_23            = 2'h0;
assign OE_DATA_123_const_net_23            = 2'h0;
assign OE_DATA_124_const_net_23            = 2'h0;
assign OE_DATA_125_const_net_23            = 2'h0;
assign OE_DATA_126_const_net_23            = 2'h0;
assign OE_DATA_127_const_net_23            = 2'h0;
assign RX_DQS_90_const_net_18              = 2'h0;
assign EYE_MONITOR_LANE_WIDTH_const_net_20 = 3'h0;
assign TX_DATA_1_const_net_19              = 8'h00;
assign TX_DATA_2_const_net_21              = 8'h00;
assign TX_DATA_3_const_net_21              = 8'h00;
assign TX_DATA_4_const_net_21              = 8'h00;
assign TX_DATA_5_const_net_21              = 8'h00;
assign TX_DATA_6_const_net_21              = 8'h00;
assign TX_DATA_7_const_net_21              = 8'h00;
assign TX_DATA_8_const_net_23              = 8'h00;
assign TX_DATA_9_const_net_23              = 8'h00;
assign TX_DATA_10_const_net_23             = 8'h00;
assign TX_DATA_11_const_net_23             = 8'h00;
assign TX_DATA_12_const_net_24             = 8'h00;
assign TX_DATA_13_const_net_24             = 8'h00;
assign TX_DATA_14_const_net_24             = 8'h00;
assign TX_DATA_15_const_net_24             = 8'h00;
assign TX_DATA_16_const_net_24             = 8'h00;
assign TX_DATA_17_const_net_24             = 8'h00;
assign TX_DATA_18_const_net_24             = 8'h00;
assign TX_DATA_19_const_net_24             = 8'h00;
assign TX_DATA_20_const_net_24             = 8'h00;
assign TX_DATA_21_const_net_24             = 8'h00;
assign TX_DATA_22_const_net_24             = 8'h00;
assign TX_DATA_23_const_net_24             = 8'h00;
assign TX_DATA_24_const_net_24             = 8'h00;
assign TX_DATA_25_const_net_24             = 8'h00;
assign TX_DATA_26_const_net_24             = 8'h00;
assign TX_DATA_27_const_net_24             = 8'h00;
assign TX_DATA_28_const_net_24             = 8'h00;
assign TX_DATA_29_const_net_24             = 8'h00;
assign TX_DATA_30_const_net_24             = 8'h00;
assign TX_DATA_31_const_net_24             = 8'h00;
assign TX_DATA_32_const_net_24             = 8'h00;
assign TX_DATA_33_const_net_24             = 8'h00;
assign TX_DATA_34_const_net_24             = 8'h00;
assign TX_DATA_35_const_net_24             = 8'h00;
assign TX_DATA_36_const_net_24             = 8'h00;
assign TX_DATA_37_const_net_24             = 8'h00;
assign TX_DATA_38_const_net_24             = 8'h00;
assign TX_DATA_39_const_net_24             = 8'h00;
assign TX_DATA_40_const_net_24             = 8'h00;
assign TX_DATA_41_const_net_24             = 8'h00;
assign TX_DATA_42_const_net_24             = 8'h00;
assign TX_DATA_43_const_net_24             = 8'h00;
assign TX_DATA_44_const_net_24             = 8'h00;
assign TX_DATA_45_const_net_24             = 8'h00;
assign TX_DATA_46_const_net_24             = 8'h00;
assign TX_DATA_47_const_net_24             = 8'h00;
assign TX_DATA_48_const_net_24             = 8'h00;
assign TX_DATA_49_const_net_24             = 8'h00;
assign TX_DATA_50_const_net_24             = 8'h00;
assign TX_DATA_51_const_net_24             = 8'h00;
assign TX_DATA_52_const_net_24             = 8'h00;
assign TX_DATA_53_const_net_24             = 8'h00;
assign TX_DATA_54_const_net_24             = 8'h00;
assign TX_DATA_55_const_net_24             = 8'h00;
assign TX_DATA_56_const_net_24             = 8'h00;
assign TX_DATA_57_const_net_24             = 8'h00;
assign TX_DATA_58_const_net_24             = 8'h00;
assign TX_DATA_59_const_net_24             = 8'h00;
assign TX_DATA_60_const_net_24             = 8'h00;
assign TX_DATA_61_const_net_24             = 8'h00;
assign TX_DATA_62_const_net_24             = 8'h00;
assign TX_DATA_63_const_net_24             = 8'h00;
assign TX_DATA_64_const_net_24             = 8'h00;
assign TX_DATA_65_const_net_24             = 8'h00;
assign TX_DATA_66_const_net_24             = 8'h00;
assign TX_DATA_67_const_net_24             = 8'h00;
assign TX_DATA_68_const_net_24             = 8'h00;
assign TX_DATA_69_const_net_24             = 8'h00;
assign TX_DATA_70_const_net_24             = 8'h00;
assign TX_DATA_71_const_net_24             = 8'h00;
assign TX_DATA_72_const_net_24             = 8'h00;
assign TX_DATA_73_const_net_24             = 8'h00;
assign TX_DATA_74_const_net_24             = 8'h00;
assign TX_DATA_75_const_net_24             = 8'h00;
assign TX_DATA_76_const_net_24             = 8'h00;
assign TX_DATA_77_const_net_24             = 8'h00;
assign TX_DATA_78_const_net_24             = 8'h00;
assign TX_DATA_79_const_net_24             = 8'h00;
assign TX_DATA_80_const_net_24             = 8'h00;
assign TX_DATA_81_const_net_24             = 8'h00;
assign TX_DATA_82_const_net_24             = 8'h00;
assign TX_DATA_83_const_net_24             = 8'h00;
assign TX_DATA_84_const_net_24             = 8'h00;
assign TX_DATA_85_const_net_24             = 8'h00;
assign TX_DATA_86_const_net_24             = 8'h00;
assign TX_DATA_87_const_net_24             = 8'h00;
assign TX_DATA_88_const_net_24             = 8'h00;
assign TX_DATA_89_const_net_24             = 8'h00;
assign TX_DATA_90_const_net_24             = 8'h00;
assign TX_DATA_91_const_net_24             = 8'h00;
assign TX_DATA_92_const_net_24             = 8'h00;
assign TX_DATA_93_const_net_24             = 8'h00;
assign TX_DATA_94_const_net_24             = 8'h00;
assign TX_DATA_95_const_net_24             = 8'h00;
assign TX_DATA_96_const_net_24             = 8'h00;
assign TX_DATA_97_const_net_24             = 8'h00;
assign TX_DATA_98_const_net_24             = 8'h00;
assign TX_DATA_99_const_net_24             = 8'h00;
assign TX_DATA_100_const_net_24            = 8'h00;
assign TX_DATA_101_const_net_24            = 8'h00;
assign TX_DATA_102_const_net_24            = 8'h00;
assign TX_DATA_103_const_net_24            = 8'h00;
assign TX_DATA_104_const_net_24            = 8'h00;
assign TX_DATA_105_const_net_24            = 8'h00;
assign TX_DATA_106_const_net_24            = 8'h00;
assign TX_DATA_107_const_net_24            = 8'h00;
assign TX_DATA_108_const_net_24            = 8'h00;
assign TX_DATA_109_const_net_24            = 8'h00;
assign TX_DATA_110_const_net_24            = 8'h00;
assign TX_DATA_111_const_net_24            = 8'h00;
assign TX_DATA_112_const_net_24            = 8'h00;
assign TX_DATA_113_const_net_24            = 8'h00;
assign TX_DATA_114_const_net_24            = 8'h00;
assign TX_DATA_115_const_net_24            = 8'h00;
assign TX_DATA_116_const_net_24            = 8'h00;
assign TX_DATA_117_const_net_24            = 8'h00;
assign TX_DATA_118_const_net_24            = 8'h00;
assign TX_DATA_119_const_net_24            = 8'h00;
assign TX_DATA_120_const_net_24            = 8'h00;
assign TX_DATA_121_const_net_24            = 8'h00;
assign TX_DATA_122_const_net_24            = 8'h00;
assign TX_DATA_123_const_net_24            = 8'h00;
assign TX_DATA_124_const_net_24            = 8'h00;
assign TX_DATA_125_const_net_24            = 8'h00;
assign TX_DATA_126_const_net_24            = 8'h00;
assign TX_DATA_127_const_net_24            = 8'h00;
assign OE_DATA_1_const_net_22              = 4'h0;
assign OE_DATA_2_const_net_22              = 4'h0;
assign OE_DATA_3_const_net_22              = 4'h0;
assign OE_DATA_4_const_net_22              = 4'h0;
assign OE_DATA_5_const_net_22              = 4'h0;
assign OE_DATA_6_const_net_22              = 4'h0;
assign OE_DATA_7_const_net_22              = 4'h0;
assign OE_DATA_8_const_net_24              = 4'h0;
assign OE_DATA_9_const_net_24              = 4'h0;
assign OE_DATA_10_const_net_24             = 4'h0;
assign OE_DATA_11_const_net_24             = 4'h0;
assign OE_DATA_12_const_net_24             = 4'h0;
assign OE_DATA_13_const_net_24             = 4'h0;
assign OE_DATA_14_const_net_24             = 4'h0;
assign OE_DATA_15_const_net_24             = 4'h0;
assign OE_DATA_16_const_net_24             = 4'h0;
assign OE_DATA_17_const_net_24             = 4'h0;
assign OE_DATA_18_const_net_24             = 4'h0;
assign OE_DATA_19_const_net_24             = 4'h0;
assign OE_DATA_20_const_net_24             = 4'h0;
assign OE_DATA_21_const_net_24             = 4'h0;
assign OE_DATA_22_const_net_24             = 4'h0;
assign OE_DATA_23_const_net_24             = 4'h0;
assign OE_DATA_24_const_net_24             = 4'h0;
assign OE_DATA_25_const_net_24             = 4'h0;
assign OE_DATA_26_const_net_24             = 4'h0;
assign OE_DATA_27_const_net_24             = 4'h0;
assign OE_DATA_28_const_net_24             = 4'h0;
assign OE_DATA_29_const_net_24             = 4'h0;
assign OE_DATA_30_const_net_24             = 4'h0;
assign OE_DATA_31_const_net_24             = 4'h0;
assign OE_DATA_32_const_net_24             = 4'h0;
assign OE_DATA_33_const_net_24             = 4'h0;
assign OE_DATA_34_const_net_24             = 4'h0;
assign OE_DATA_35_const_net_24             = 4'h0;
assign OE_DATA_36_const_net_24             = 4'h0;
assign OE_DATA_37_const_net_24             = 4'h0;
assign OE_DATA_38_const_net_24             = 4'h0;
assign OE_DATA_39_const_net_24             = 4'h0;
assign OE_DATA_40_const_net_24             = 4'h0;
assign OE_DATA_41_const_net_24             = 4'h0;
assign OE_DATA_42_const_net_24             = 4'h0;
assign OE_DATA_43_const_net_24             = 4'h0;
assign OE_DATA_44_const_net_24             = 4'h0;
assign OE_DATA_45_const_net_24             = 4'h0;
assign OE_DATA_46_const_net_24             = 4'h0;
assign OE_DATA_47_const_net_24             = 4'h0;
assign OE_DATA_48_const_net_24             = 4'h0;
assign OE_DATA_49_const_net_24             = 4'h0;
assign OE_DATA_50_const_net_24             = 4'h0;
assign OE_DATA_51_const_net_24             = 4'h0;
assign OE_DATA_52_const_net_24             = 4'h0;
assign OE_DATA_53_const_net_24             = 4'h0;
assign OE_DATA_54_const_net_24             = 4'h0;
assign OE_DATA_55_const_net_24             = 4'h0;
assign OE_DATA_56_const_net_24             = 4'h0;
assign OE_DATA_57_const_net_24             = 4'h0;
assign OE_DATA_58_const_net_24             = 4'h0;
assign OE_DATA_59_const_net_24             = 4'h0;
assign OE_DATA_60_const_net_24             = 4'h0;
assign OE_DATA_61_const_net_24             = 4'h0;
assign OE_DATA_62_const_net_24             = 4'h0;
assign OE_DATA_63_const_net_24             = 4'h0;
assign OE_DATA_64_const_net_24             = 4'h0;
assign OE_DATA_65_const_net_24             = 4'h0;
assign OE_DATA_66_const_net_24             = 4'h0;
assign OE_DATA_67_const_net_24             = 4'h0;
assign OE_DATA_68_const_net_24             = 4'h0;
assign OE_DATA_69_const_net_24             = 4'h0;
assign OE_DATA_70_const_net_24             = 4'h0;
assign OE_DATA_71_const_net_24             = 4'h0;
assign OE_DATA_72_const_net_24             = 4'h0;
assign OE_DATA_73_const_net_24             = 4'h0;
assign OE_DATA_74_const_net_24             = 4'h0;
assign OE_DATA_75_const_net_24             = 4'h0;
assign OE_DATA_76_const_net_24             = 4'h0;
assign OE_DATA_77_const_net_24             = 4'h0;
assign OE_DATA_78_const_net_24             = 4'h0;
assign OE_DATA_79_const_net_24             = 4'h0;
assign OE_DATA_80_const_net_24             = 4'h0;
assign OE_DATA_81_const_net_24             = 4'h0;
assign OE_DATA_82_const_net_24             = 4'h0;
assign OE_DATA_83_const_net_24             = 4'h0;
assign OE_DATA_84_const_net_24             = 4'h0;
assign OE_DATA_85_const_net_24             = 4'h0;
assign OE_DATA_86_const_net_24             = 4'h0;
assign OE_DATA_87_const_net_24             = 4'h0;
assign OE_DATA_88_const_net_24             = 4'h0;
assign OE_DATA_89_const_net_24             = 4'h0;
assign OE_DATA_90_const_net_24             = 4'h0;
assign OE_DATA_91_const_net_24             = 4'h0;
assign OE_DATA_92_const_net_24             = 4'h0;
assign OE_DATA_93_const_net_24             = 4'h0;
assign OE_DATA_94_const_net_24             = 4'h0;
assign OE_DATA_95_const_net_24             = 4'h0;
assign OE_DATA_96_const_net_24             = 4'h0;
assign OE_DATA_97_const_net_24             = 4'h0;
assign OE_DATA_98_const_net_24             = 4'h0;
assign OE_DATA_99_const_net_24             = 4'h0;
assign OE_DATA_100_const_net_24            = 4'h0;
assign OE_DATA_101_const_net_24            = 4'h0;
assign OE_DATA_102_const_net_24            = 4'h0;
assign OE_DATA_103_const_net_24            = 4'h0;
assign OE_DATA_104_const_net_24            = 4'h0;
assign OE_DATA_105_const_net_24            = 4'h0;
assign OE_DATA_106_const_net_24            = 4'h0;
assign OE_DATA_107_const_net_24            = 4'h0;
assign OE_DATA_108_const_net_24            = 4'h0;
assign OE_DATA_109_const_net_24            = 4'h0;
assign OE_DATA_110_const_net_24            = 4'h0;
assign OE_DATA_111_const_net_24            = 4'h0;
assign OE_DATA_112_const_net_24            = 4'h0;
assign OE_DATA_113_const_net_24            = 4'h0;
assign OE_DATA_114_const_net_24            = 4'h0;
assign OE_DATA_115_const_net_24            = 4'h0;
assign OE_DATA_116_const_net_24            = 4'h0;
assign OE_DATA_117_const_net_24            = 4'h0;
assign OE_DATA_118_const_net_24            = 4'h0;
assign OE_DATA_119_const_net_24            = 4'h0;
assign OE_DATA_120_const_net_24            = 4'h0;
assign OE_DATA_121_const_net_24            = 4'h0;
assign OE_DATA_122_const_net_24            = 4'h0;
assign OE_DATA_123_const_net_24            = 4'h0;
assign OE_DATA_124_const_net_24            = 4'h0;
assign OE_DATA_125_const_net_24            = 4'h0;
assign OE_DATA_126_const_net_24            = 4'h0;
assign OE_DATA_127_const_net_24            = 4'h0;
assign CDR_CLK_B_SEL_const_net_2           = 11'h000;
assign FIFO_WR_PTR_const_net_19            = 3'h0;
assign FIFO_RD_PTR_const_net_19            = 3'h0;
assign EYE_MONITOR_LANE_WIDTH_const_net_21 = 3'h0;
assign TX_DATA_1_const_net_20              = 8'h00;
assign TX_DATA_2_const_net_22              = 8'h00;
assign TX_DATA_3_const_net_22              = 8'h00;
assign TX_DATA_4_const_net_22              = 8'h00;
assign TX_DATA_5_const_net_22              = 8'h00;
assign TX_DATA_6_const_net_22              = 8'h00;
assign TX_DATA_7_const_net_22              = 8'h00;
assign TX_DATA_8_const_net_24              = 8'h00;
assign TX_DATA_9_const_net_24              = 8'h00;
assign TX_DATA_10_const_net_24             = 8'h00;
assign TX_DATA_11_const_net_24             = 8'h00;
assign TX_DATA_12_const_net_25             = 8'h00;
assign TX_DATA_13_const_net_25             = 8'h00;
assign TX_DATA_14_const_net_25             = 8'h00;
assign TX_DATA_15_const_net_25             = 8'h00;
assign TX_DATA_16_const_net_25             = 8'h00;
assign TX_DATA_17_const_net_25             = 8'h00;
assign TX_DATA_18_const_net_25             = 8'h00;
assign TX_DATA_19_const_net_25             = 8'h00;
assign TX_DATA_20_const_net_25             = 8'h00;
assign TX_DATA_21_const_net_25             = 8'h00;
assign TX_DATA_22_const_net_25             = 8'h00;
assign TX_DATA_23_const_net_25             = 8'h00;
assign TX_DATA_24_const_net_25             = 8'h00;
assign TX_DATA_25_const_net_25             = 8'h00;
assign TX_DATA_26_const_net_25             = 8'h00;
assign TX_DATA_27_const_net_25             = 8'h00;
assign TX_DATA_28_const_net_25             = 8'h00;
assign TX_DATA_29_const_net_25             = 8'h00;
assign TX_DATA_30_const_net_25             = 8'h00;
assign TX_DATA_31_const_net_25             = 8'h00;
assign TX_DATA_32_const_net_25             = 8'h00;
assign TX_DATA_33_const_net_25             = 8'h00;
assign TX_DATA_34_const_net_25             = 8'h00;
assign TX_DATA_35_const_net_25             = 8'h00;
assign TX_DATA_36_const_net_25             = 8'h00;
assign TX_DATA_37_const_net_25             = 8'h00;
assign TX_DATA_38_const_net_25             = 8'h00;
assign TX_DATA_39_const_net_25             = 8'h00;
assign TX_DATA_40_const_net_25             = 8'h00;
assign TX_DATA_41_const_net_25             = 8'h00;
assign TX_DATA_42_const_net_25             = 8'h00;
assign TX_DATA_43_const_net_25             = 8'h00;
assign TX_DATA_44_const_net_25             = 8'h00;
assign TX_DATA_45_const_net_25             = 8'h00;
assign TX_DATA_46_const_net_25             = 8'h00;
assign TX_DATA_47_const_net_25             = 8'h00;
assign TX_DATA_48_const_net_25             = 8'h00;
assign TX_DATA_49_const_net_25             = 8'h00;
assign TX_DATA_50_const_net_25             = 8'h00;
assign TX_DATA_51_const_net_25             = 8'h00;
assign TX_DATA_52_const_net_25             = 8'h00;
assign TX_DATA_53_const_net_25             = 8'h00;
assign TX_DATA_54_const_net_25             = 8'h00;
assign TX_DATA_55_const_net_25             = 8'h00;
assign TX_DATA_56_const_net_25             = 8'h00;
assign TX_DATA_57_const_net_25             = 8'h00;
assign TX_DATA_58_const_net_25             = 8'h00;
assign TX_DATA_59_const_net_25             = 8'h00;
assign TX_DATA_60_const_net_25             = 8'h00;
assign TX_DATA_61_const_net_25             = 8'h00;
assign TX_DATA_62_const_net_25             = 8'h00;
assign TX_DATA_63_const_net_25             = 8'h00;
assign TX_DATA_64_const_net_25             = 8'h00;
assign TX_DATA_65_const_net_25             = 8'h00;
assign TX_DATA_66_const_net_25             = 8'h00;
assign TX_DATA_67_const_net_25             = 8'h00;
assign TX_DATA_68_const_net_25             = 8'h00;
assign TX_DATA_69_const_net_25             = 8'h00;
assign TX_DATA_70_const_net_25             = 8'h00;
assign TX_DATA_71_const_net_25             = 8'h00;
assign TX_DATA_72_const_net_25             = 8'h00;
assign TX_DATA_73_const_net_25             = 8'h00;
assign TX_DATA_74_const_net_25             = 8'h00;
assign TX_DATA_75_const_net_25             = 8'h00;
assign TX_DATA_76_const_net_25             = 8'h00;
assign TX_DATA_77_const_net_25             = 8'h00;
assign TX_DATA_78_const_net_25             = 8'h00;
assign TX_DATA_79_const_net_25             = 8'h00;
assign TX_DATA_80_const_net_25             = 8'h00;
assign TX_DATA_81_const_net_25             = 8'h00;
assign TX_DATA_82_const_net_25             = 8'h00;
assign TX_DATA_83_const_net_25             = 8'h00;
assign TX_DATA_84_const_net_25             = 8'h00;
assign TX_DATA_85_const_net_25             = 8'h00;
assign TX_DATA_86_const_net_25             = 8'h00;
assign TX_DATA_87_const_net_25             = 8'h00;
assign TX_DATA_88_const_net_25             = 8'h00;
assign TX_DATA_89_const_net_25             = 8'h00;
assign TX_DATA_90_const_net_25             = 8'h00;
assign TX_DATA_91_const_net_25             = 8'h00;
assign TX_DATA_92_const_net_25             = 8'h00;
assign TX_DATA_93_const_net_25             = 8'h00;
assign TX_DATA_94_const_net_25             = 8'h00;
assign TX_DATA_95_const_net_25             = 8'h00;
assign TX_DATA_96_const_net_25             = 8'h00;
assign TX_DATA_97_const_net_25             = 8'h00;
assign TX_DATA_98_const_net_25             = 8'h00;
assign TX_DATA_99_const_net_25             = 8'h00;
assign TX_DATA_100_const_net_25            = 8'h00;
assign TX_DATA_101_const_net_25            = 8'h00;
assign TX_DATA_102_const_net_25            = 8'h00;
assign TX_DATA_103_const_net_25            = 8'h00;
assign TX_DATA_104_const_net_25            = 8'h00;
assign TX_DATA_105_const_net_25            = 8'h00;
assign TX_DATA_106_const_net_25            = 8'h00;
assign TX_DATA_107_const_net_25            = 8'h00;
assign TX_DATA_108_const_net_25            = 8'h00;
assign TX_DATA_109_const_net_25            = 8'h00;
assign TX_DATA_110_const_net_25            = 8'h00;
assign TX_DATA_111_const_net_25            = 8'h00;
assign TX_DATA_112_const_net_25            = 8'h00;
assign TX_DATA_113_const_net_25            = 8'h00;
assign TX_DATA_114_const_net_25            = 8'h00;
assign TX_DATA_115_const_net_25            = 8'h00;
assign TX_DATA_116_const_net_25            = 8'h00;
assign TX_DATA_117_const_net_25            = 8'h00;
assign TX_DATA_118_const_net_25            = 8'h00;
assign TX_DATA_119_const_net_25            = 8'h00;
assign TX_DATA_120_const_net_25            = 8'h00;
assign TX_DATA_121_const_net_25            = 8'h00;
assign TX_DATA_122_const_net_25            = 8'h00;
assign TX_DATA_123_const_net_25            = 8'h00;
assign TX_DATA_124_const_net_25            = 8'h00;
assign TX_DATA_125_const_net_25            = 8'h00;
assign TX_DATA_126_const_net_25            = 8'h00;
assign TX_DATA_127_const_net_25            = 8'h00;
assign OE_DATA_1_const_net_23              = 4'h0;
assign OE_DATA_2_const_net_23              = 4'h0;
assign OE_DATA_3_const_net_23              = 4'h0;
assign OE_DATA_4_const_net_23              = 4'h0;
assign OE_DATA_5_const_net_23              = 4'h0;
assign OE_DATA_6_const_net_23              = 4'h0;
assign OE_DATA_7_const_net_23              = 4'h0;
assign OE_DATA_8_const_net_25              = 4'h0;
assign OE_DATA_9_const_net_25              = 4'h0;
assign OE_DATA_10_const_net_25             = 4'h0;
assign OE_DATA_11_const_net_25             = 4'h0;
assign OE_DATA_12_const_net_25             = 4'h0;
assign OE_DATA_13_const_net_25             = 4'h0;
assign OE_DATA_14_const_net_25             = 4'h0;
assign OE_DATA_15_const_net_25             = 4'h0;
assign OE_DATA_16_const_net_25             = 4'h0;
assign OE_DATA_17_const_net_25             = 4'h0;
assign OE_DATA_18_const_net_25             = 4'h0;
assign OE_DATA_19_const_net_25             = 4'h0;
assign OE_DATA_20_const_net_25             = 4'h0;
assign OE_DATA_21_const_net_25             = 4'h0;
assign OE_DATA_22_const_net_25             = 4'h0;
assign OE_DATA_23_const_net_25             = 4'h0;
assign OE_DATA_24_const_net_25             = 4'h0;
assign OE_DATA_25_const_net_25             = 4'h0;
assign OE_DATA_26_const_net_25             = 4'h0;
assign OE_DATA_27_const_net_25             = 4'h0;
assign OE_DATA_28_const_net_25             = 4'h0;
assign OE_DATA_29_const_net_25             = 4'h0;
assign OE_DATA_30_const_net_25             = 4'h0;
assign OE_DATA_31_const_net_25             = 4'h0;
assign OE_DATA_32_const_net_25             = 4'h0;
assign OE_DATA_33_const_net_25             = 4'h0;
assign OE_DATA_34_const_net_25             = 4'h0;
assign OE_DATA_35_const_net_25             = 4'h0;
assign OE_DATA_36_const_net_25             = 4'h0;
assign OE_DATA_37_const_net_25             = 4'h0;
assign OE_DATA_38_const_net_25             = 4'h0;
assign OE_DATA_39_const_net_25             = 4'h0;
assign OE_DATA_40_const_net_25             = 4'h0;
assign OE_DATA_41_const_net_25             = 4'h0;
assign OE_DATA_42_const_net_25             = 4'h0;
assign OE_DATA_43_const_net_25             = 4'h0;
assign OE_DATA_44_const_net_25             = 4'h0;
assign OE_DATA_45_const_net_25             = 4'h0;
assign OE_DATA_46_const_net_25             = 4'h0;
assign OE_DATA_47_const_net_25             = 4'h0;
assign OE_DATA_48_const_net_25             = 4'h0;
assign OE_DATA_49_const_net_25             = 4'h0;
assign OE_DATA_50_const_net_25             = 4'h0;
assign OE_DATA_51_const_net_25             = 4'h0;
assign OE_DATA_52_const_net_25             = 4'h0;
assign OE_DATA_53_const_net_25             = 4'h0;
assign OE_DATA_54_const_net_25             = 4'h0;
assign OE_DATA_55_const_net_25             = 4'h0;
assign OE_DATA_56_const_net_25             = 4'h0;
assign OE_DATA_57_const_net_25             = 4'h0;
assign OE_DATA_58_const_net_25             = 4'h0;
assign OE_DATA_59_const_net_25             = 4'h0;
assign OE_DATA_60_const_net_25             = 4'h0;
assign OE_DATA_61_const_net_25             = 4'h0;
assign OE_DATA_62_const_net_25             = 4'h0;
assign OE_DATA_63_const_net_25             = 4'h0;
assign OE_DATA_64_const_net_25             = 4'h0;
assign OE_DATA_65_const_net_25             = 4'h0;
assign OE_DATA_66_const_net_25             = 4'h0;
assign OE_DATA_67_const_net_25             = 4'h0;
assign OE_DATA_68_const_net_25             = 4'h0;
assign OE_DATA_69_const_net_25             = 4'h0;
assign OE_DATA_70_const_net_25             = 4'h0;
assign OE_DATA_71_const_net_25             = 4'h0;
assign OE_DATA_72_const_net_25             = 4'h0;
assign OE_DATA_73_const_net_25             = 4'h0;
assign OE_DATA_74_const_net_25             = 4'h0;
assign OE_DATA_75_const_net_25             = 4'h0;
assign OE_DATA_76_const_net_25             = 4'h0;
assign OE_DATA_77_const_net_25             = 4'h0;
assign OE_DATA_78_const_net_25             = 4'h0;
assign OE_DATA_79_const_net_25             = 4'h0;
assign OE_DATA_80_const_net_25             = 4'h0;
assign OE_DATA_81_const_net_25             = 4'h0;
assign OE_DATA_82_const_net_25             = 4'h0;
assign OE_DATA_83_const_net_25             = 4'h0;
assign OE_DATA_84_const_net_25             = 4'h0;
assign OE_DATA_85_const_net_25             = 4'h0;
assign OE_DATA_86_const_net_25             = 4'h0;
assign OE_DATA_87_const_net_25             = 4'h0;
assign OE_DATA_88_const_net_25             = 4'h0;
assign OE_DATA_89_const_net_25             = 4'h0;
assign OE_DATA_90_const_net_25             = 4'h0;
assign OE_DATA_91_const_net_25             = 4'h0;
assign OE_DATA_92_const_net_25             = 4'h0;
assign OE_DATA_93_const_net_25             = 4'h0;
assign OE_DATA_94_const_net_25             = 4'h0;
assign OE_DATA_95_const_net_25             = 4'h0;
assign OE_DATA_96_const_net_25             = 4'h0;
assign OE_DATA_97_const_net_25             = 4'h0;
assign OE_DATA_98_const_net_25             = 4'h0;
assign OE_DATA_99_const_net_25             = 4'h0;
assign OE_DATA_100_const_net_25            = 4'h0;
assign OE_DATA_101_const_net_25            = 4'h0;
assign OE_DATA_102_const_net_25            = 4'h0;
assign OE_DATA_103_const_net_25            = 4'h0;
assign OE_DATA_104_const_net_25            = 4'h0;
assign OE_DATA_105_const_net_25            = 4'h0;
assign OE_DATA_106_const_net_25            = 4'h0;
assign OE_DATA_107_const_net_25            = 4'h0;
assign OE_DATA_108_const_net_25            = 4'h0;
assign OE_DATA_109_const_net_25            = 4'h0;
assign OE_DATA_110_const_net_25            = 4'h0;
assign OE_DATA_111_const_net_25            = 4'h0;
assign OE_DATA_112_const_net_25            = 4'h0;
assign OE_DATA_113_const_net_25            = 4'h0;
assign OE_DATA_114_const_net_25            = 4'h0;
assign OE_DATA_115_const_net_25            = 4'h0;
assign OE_DATA_116_const_net_25            = 4'h0;
assign OE_DATA_117_const_net_25            = 4'h0;
assign OE_DATA_118_const_net_25            = 4'h0;
assign OE_DATA_119_const_net_25            = 4'h0;
assign OE_DATA_120_const_net_25            = 4'h0;
assign OE_DATA_121_const_net_25            = 4'h0;
assign OE_DATA_122_const_net_25            = 4'h0;
assign OE_DATA_123_const_net_25            = 4'h0;
assign OE_DATA_124_const_net_25            = 4'h0;
assign OE_DATA_125_const_net_25            = 4'h0;
assign OE_DATA_126_const_net_25            = 4'h0;
assign OE_DATA_127_const_net_25            = 4'h0;
assign TX_DATA_8_const_net_25              = 8'h00;
assign TX_DATA_9_const_net_25              = 8'h00;
assign TX_DATA_10_const_net_25             = 8'h00;
assign TX_DATA_11_const_net_25             = 8'h00;
assign TX_DATA_12_const_net_26             = 8'h00;
assign TX_DATA_13_const_net_26             = 8'h00;
assign TX_DATA_14_const_net_26             = 8'h00;
assign TX_DATA_15_const_net_26             = 8'h00;
assign TX_DATA_16_const_net_26             = 8'h00;
assign TX_DATA_17_const_net_26             = 8'h00;
assign TX_DATA_18_const_net_26             = 8'h00;
assign TX_DATA_19_const_net_26             = 8'h00;
assign TX_DATA_20_const_net_26             = 8'h00;
assign TX_DATA_21_const_net_26             = 8'h00;
assign TX_DATA_22_const_net_26             = 8'h00;
assign TX_DATA_23_const_net_26             = 8'h00;
assign TX_DATA_24_const_net_26             = 8'h00;
assign TX_DATA_25_const_net_26             = 8'h00;
assign TX_DATA_26_const_net_26             = 8'h00;
assign TX_DATA_27_const_net_26             = 8'h00;
assign TX_DATA_28_const_net_26             = 8'h00;
assign TX_DATA_29_const_net_26             = 8'h00;
assign TX_DATA_30_const_net_26             = 8'h00;
assign TX_DATA_31_const_net_26             = 8'h00;
assign TX_DATA_32_const_net_26             = 8'h00;
assign TX_DATA_33_const_net_26             = 8'h00;
assign TX_DATA_34_const_net_26             = 8'h00;
assign TX_DATA_35_const_net_26             = 8'h00;
assign TX_DATA_36_const_net_26             = 8'h00;
assign TX_DATA_37_const_net_26             = 8'h00;
assign TX_DATA_38_const_net_26             = 8'h00;
assign TX_DATA_39_const_net_26             = 8'h00;
assign TX_DATA_40_const_net_26             = 8'h00;
assign TX_DATA_41_const_net_26             = 8'h00;
assign TX_DATA_42_const_net_26             = 8'h00;
assign TX_DATA_43_const_net_26             = 8'h00;
assign TX_DATA_44_const_net_26             = 8'h00;
assign TX_DATA_45_const_net_26             = 8'h00;
assign TX_DATA_46_const_net_26             = 8'h00;
assign TX_DATA_47_const_net_26             = 8'h00;
assign TX_DATA_48_const_net_26             = 8'h00;
assign TX_DATA_49_const_net_26             = 8'h00;
assign TX_DATA_50_const_net_26             = 8'h00;
assign TX_DATA_51_const_net_26             = 8'h00;
assign TX_DATA_52_const_net_26             = 8'h00;
assign TX_DATA_53_const_net_26             = 8'h00;
assign TX_DATA_54_const_net_26             = 8'h00;
assign TX_DATA_55_const_net_26             = 8'h00;
assign TX_DATA_56_const_net_26             = 8'h00;
assign TX_DATA_57_const_net_26             = 8'h00;
assign TX_DATA_58_const_net_26             = 8'h00;
assign TX_DATA_59_const_net_26             = 8'h00;
assign TX_DATA_60_const_net_26             = 8'h00;
assign TX_DATA_61_const_net_26             = 8'h00;
assign TX_DATA_62_const_net_26             = 8'h00;
assign TX_DATA_63_const_net_26             = 8'h00;
assign TX_DATA_64_const_net_26             = 8'h00;
assign TX_DATA_65_const_net_26             = 8'h00;
assign TX_DATA_66_const_net_26             = 8'h00;
assign TX_DATA_67_const_net_26             = 8'h00;
assign TX_DATA_68_const_net_26             = 8'h00;
assign TX_DATA_69_const_net_26             = 8'h00;
assign TX_DATA_70_const_net_26             = 8'h00;
assign TX_DATA_71_const_net_26             = 8'h00;
assign TX_DATA_72_const_net_26             = 8'h00;
assign TX_DATA_73_const_net_26             = 8'h00;
assign TX_DATA_74_const_net_26             = 8'h00;
assign TX_DATA_75_const_net_26             = 8'h00;
assign TX_DATA_76_const_net_26             = 8'h00;
assign TX_DATA_77_const_net_26             = 8'h00;
assign TX_DATA_78_const_net_26             = 8'h00;
assign TX_DATA_79_const_net_26             = 8'h00;
assign TX_DATA_80_const_net_26             = 8'h00;
assign TX_DATA_81_const_net_26             = 8'h00;
assign TX_DATA_82_const_net_26             = 8'h00;
assign TX_DATA_83_const_net_26             = 8'h00;
assign TX_DATA_84_const_net_26             = 8'h00;
assign TX_DATA_85_const_net_26             = 8'h00;
assign TX_DATA_86_const_net_26             = 8'h00;
assign TX_DATA_87_const_net_26             = 8'h00;
assign TX_DATA_88_const_net_26             = 8'h00;
assign TX_DATA_89_const_net_26             = 8'h00;
assign TX_DATA_90_const_net_26             = 8'h00;
assign TX_DATA_91_const_net_26             = 8'h00;
assign TX_DATA_92_const_net_26             = 8'h00;
assign TX_DATA_93_const_net_26             = 8'h00;
assign TX_DATA_94_const_net_26             = 8'h00;
assign TX_DATA_95_const_net_26             = 8'h00;
assign TX_DATA_96_const_net_26             = 8'h00;
assign TX_DATA_97_const_net_26             = 8'h00;
assign TX_DATA_98_const_net_26             = 8'h00;
assign TX_DATA_99_const_net_26             = 8'h00;
assign TX_DATA_100_const_net_26            = 8'h00;
assign TX_DATA_101_const_net_26            = 8'h00;
assign TX_DATA_102_const_net_26            = 8'h00;
assign TX_DATA_103_const_net_26            = 8'h00;
assign TX_DATA_104_const_net_26            = 8'h00;
assign TX_DATA_105_const_net_26            = 8'h00;
assign TX_DATA_106_const_net_26            = 8'h00;
assign TX_DATA_107_const_net_26            = 8'h00;
assign TX_DATA_108_const_net_26            = 8'h00;
assign TX_DATA_109_const_net_26            = 8'h00;
assign TX_DATA_110_const_net_26            = 8'h00;
assign TX_DATA_111_const_net_26            = 8'h00;
assign TX_DATA_112_const_net_26            = 8'h00;
assign TX_DATA_113_const_net_26            = 8'h00;
assign TX_DATA_114_const_net_26            = 8'h00;
assign TX_DATA_115_const_net_26            = 8'h00;
assign TX_DATA_116_const_net_26            = 8'h00;
assign TX_DATA_117_const_net_26            = 8'h00;
assign TX_DATA_118_const_net_26            = 8'h00;
assign TX_DATA_119_const_net_26            = 8'h00;
assign TX_DATA_120_const_net_26            = 8'h00;
assign TX_DATA_121_const_net_26            = 8'h00;
assign TX_DATA_122_const_net_26            = 8'h00;
assign TX_DATA_123_const_net_26            = 8'h00;
assign TX_DATA_124_const_net_26            = 8'h00;
assign TX_DATA_125_const_net_26            = 8'h00;
assign TX_DATA_126_const_net_26            = 8'h00;
assign TX_DATA_127_const_net_26            = 8'h00;
assign OE_DATA_8_const_net_26              = 4'h0;
assign OE_DATA_9_const_net_26              = 4'h0;
assign OE_DATA_10_const_net_26             = 4'h0;
assign OE_DATA_11_const_net_26             = 4'h0;
assign OE_DATA_12_const_net_26             = 4'h0;
assign OE_DATA_13_const_net_26             = 4'h0;
assign OE_DATA_14_const_net_26             = 4'h0;
assign OE_DATA_15_const_net_26             = 4'h0;
assign OE_DATA_16_const_net_26             = 4'h0;
assign OE_DATA_17_const_net_26             = 4'h0;
assign OE_DATA_18_const_net_26             = 4'h0;
assign OE_DATA_19_const_net_26             = 4'h0;
assign OE_DATA_20_const_net_26             = 4'h0;
assign OE_DATA_21_const_net_26             = 4'h0;
assign OE_DATA_22_const_net_26             = 4'h0;
assign OE_DATA_23_const_net_26             = 4'h0;
assign OE_DATA_24_const_net_26             = 4'h0;
assign OE_DATA_25_const_net_26             = 4'h0;
assign OE_DATA_26_const_net_26             = 4'h0;
assign OE_DATA_27_const_net_26             = 4'h0;
assign OE_DATA_28_const_net_26             = 4'h0;
assign OE_DATA_29_const_net_26             = 4'h0;
assign OE_DATA_30_const_net_26             = 4'h0;
assign OE_DATA_31_const_net_26             = 4'h0;
assign OE_DATA_32_const_net_26             = 4'h0;
assign OE_DATA_33_const_net_26             = 4'h0;
assign OE_DATA_34_const_net_26             = 4'h0;
assign OE_DATA_35_const_net_26             = 4'h0;
assign OE_DATA_36_const_net_26             = 4'h0;
assign OE_DATA_37_const_net_26             = 4'h0;
assign OE_DATA_38_const_net_26             = 4'h0;
assign OE_DATA_39_const_net_26             = 4'h0;
assign OE_DATA_40_const_net_26             = 4'h0;
assign OE_DATA_41_const_net_26             = 4'h0;
assign OE_DATA_42_const_net_26             = 4'h0;
assign OE_DATA_43_const_net_26             = 4'h0;
assign OE_DATA_44_const_net_26             = 4'h0;
assign OE_DATA_45_const_net_26             = 4'h0;
assign OE_DATA_46_const_net_26             = 4'h0;
assign OE_DATA_47_const_net_26             = 4'h0;
assign OE_DATA_48_const_net_26             = 4'h0;
assign OE_DATA_49_const_net_26             = 4'h0;
assign OE_DATA_50_const_net_26             = 4'h0;
assign OE_DATA_51_const_net_26             = 4'h0;
assign OE_DATA_52_const_net_26             = 4'h0;
assign OE_DATA_53_const_net_26             = 4'h0;
assign OE_DATA_54_const_net_26             = 4'h0;
assign OE_DATA_55_const_net_26             = 4'h0;
assign OE_DATA_56_const_net_26             = 4'h0;
assign OE_DATA_57_const_net_26             = 4'h0;
assign OE_DATA_58_const_net_26             = 4'h0;
assign OE_DATA_59_const_net_26             = 4'h0;
assign OE_DATA_60_const_net_26             = 4'h0;
assign OE_DATA_61_const_net_26             = 4'h0;
assign OE_DATA_62_const_net_26             = 4'h0;
assign OE_DATA_63_const_net_26             = 4'h0;
assign OE_DATA_64_const_net_26             = 4'h0;
assign OE_DATA_65_const_net_26             = 4'h0;
assign OE_DATA_66_const_net_26             = 4'h0;
assign OE_DATA_67_const_net_26             = 4'h0;
assign OE_DATA_68_const_net_26             = 4'h0;
assign OE_DATA_69_const_net_26             = 4'h0;
assign OE_DATA_70_const_net_26             = 4'h0;
assign OE_DATA_71_const_net_26             = 4'h0;
assign OE_DATA_72_const_net_26             = 4'h0;
assign OE_DATA_73_const_net_26             = 4'h0;
assign OE_DATA_74_const_net_26             = 4'h0;
assign OE_DATA_75_const_net_26             = 4'h0;
assign OE_DATA_76_const_net_26             = 4'h0;
assign OE_DATA_77_const_net_26             = 4'h0;
assign OE_DATA_78_const_net_26             = 4'h0;
assign OE_DATA_79_const_net_26             = 4'h0;
assign OE_DATA_80_const_net_26             = 4'h0;
assign OE_DATA_81_const_net_26             = 4'h0;
assign OE_DATA_82_const_net_26             = 4'h0;
assign OE_DATA_83_const_net_26             = 4'h0;
assign OE_DATA_84_const_net_26             = 4'h0;
assign OE_DATA_85_const_net_26             = 4'h0;
assign OE_DATA_86_const_net_26             = 4'h0;
assign OE_DATA_87_const_net_26             = 4'h0;
assign OE_DATA_88_const_net_26             = 4'h0;
assign OE_DATA_89_const_net_26             = 4'h0;
assign OE_DATA_90_const_net_26             = 4'h0;
assign OE_DATA_91_const_net_26             = 4'h0;
assign OE_DATA_92_const_net_26             = 4'h0;
assign OE_DATA_93_const_net_26             = 4'h0;
assign OE_DATA_94_const_net_26             = 4'h0;
assign OE_DATA_95_const_net_26             = 4'h0;
assign OE_DATA_96_const_net_26             = 4'h0;
assign OE_DATA_97_const_net_26             = 4'h0;
assign OE_DATA_98_const_net_26             = 4'h0;
assign OE_DATA_99_const_net_26             = 4'h0;
assign OE_DATA_100_const_net_26            = 4'h0;
assign OE_DATA_101_const_net_26            = 4'h0;
assign OE_DATA_102_const_net_26            = 4'h0;
assign OE_DATA_103_const_net_26            = 4'h0;
assign OE_DATA_104_const_net_26            = 4'h0;
assign OE_DATA_105_const_net_26            = 4'h0;
assign OE_DATA_106_const_net_26            = 4'h0;
assign OE_DATA_107_const_net_26            = 4'h0;
assign OE_DATA_108_const_net_26            = 4'h0;
assign OE_DATA_109_const_net_26            = 4'h0;
assign OE_DATA_110_const_net_26            = 4'h0;
assign OE_DATA_111_const_net_26            = 4'h0;
assign OE_DATA_112_const_net_26            = 4'h0;
assign OE_DATA_113_const_net_26            = 4'h0;
assign OE_DATA_114_const_net_26            = 4'h0;
assign OE_DATA_115_const_net_26            = 4'h0;
assign OE_DATA_116_const_net_26            = 4'h0;
assign OE_DATA_117_const_net_26            = 4'h0;
assign OE_DATA_118_const_net_26            = 4'h0;
assign OE_DATA_119_const_net_26            = 4'h0;
assign OE_DATA_120_const_net_26            = 4'h0;
assign OE_DATA_121_const_net_26            = 4'h0;
assign OE_DATA_122_const_net_26            = 4'h0;
assign OE_DATA_123_const_net_26            = 4'h0;
assign OE_DATA_124_const_net_26            = 4'h0;
assign OE_DATA_125_const_net_26            = 4'h0;
assign OE_DATA_126_const_net_26            = 4'h0;
assign OE_DATA_127_const_net_26            = 4'h0;
assign PAD_I_const_net_5                   = 8'h00;
assign PAD_N_const_net_5                   = 8'h00;
assign PAD_I_N_const_net_5                 = 8'h00;
assign TX_DATA_1_const_net_21              = 8'h00;
assign TX_DATA_2_const_net_23              = 8'h00;
assign TX_DATA_3_const_net_23              = 8'h00;
assign TX_DATA_4_const_net_23              = 8'h00;
assign TX_DATA_5_const_net_23              = 8'h00;
assign TX_DATA_6_const_net_23              = 8'h00;
assign TX_DATA_7_const_net_23              = 8'h00;
assign TX_DATA_8_const_net_26              = 8'h00;
assign TX_DATA_9_const_net_26              = 8'h00;
assign TX_DATA_10_const_net_26             = 8'h00;
assign TX_DATA_11_const_net_26             = 8'h00;
assign TX_DATA_12_const_net_27             = 8'h00;
assign TX_DATA_13_const_net_27             = 8'h00;
assign TX_DATA_14_const_net_27             = 8'h00;
assign TX_DATA_15_const_net_27             = 8'h00;
assign TX_DATA_16_const_net_27             = 8'h00;
assign TX_DATA_17_const_net_27             = 8'h00;
assign TX_DATA_18_const_net_27             = 8'h00;
assign TX_DATA_19_const_net_27             = 8'h00;
assign TX_DATA_20_const_net_27             = 8'h00;
assign TX_DATA_21_const_net_27             = 8'h00;
assign TX_DATA_22_const_net_27             = 8'h00;
assign TX_DATA_23_const_net_27             = 8'h00;
assign TX_DATA_24_const_net_27             = 8'h00;
assign TX_DATA_25_const_net_27             = 8'h00;
assign TX_DATA_26_const_net_27             = 8'h00;
assign TX_DATA_27_const_net_27             = 8'h00;
assign TX_DATA_28_const_net_27             = 8'h00;
assign TX_DATA_29_const_net_27             = 8'h00;
assign TX_DATA_30_const_net_27             = 8'h00;
assign TX_DATA_31_const_net_27             = 8'h00;
assign TX_DATA_32_const_net_27             = 8'h00;
assign TX_DATA_33_const_net_27             = 8'h00;
assign TX_DATA_34_const_net_27             = 8'h00;
assign TX_DATA_35_const_net_27             = 8'h00;
assign TX_DATA_36_const_net_27             = 8'h00;
assign TX_DATA_37_const_net_27             = 8'h00;
assign TX_DATA_38_const_net_27             = 8'h00;
assign TX_DATA_39_const_net_27             = 8'h00;
assign TX_DATA_40_const_net_27             = 8'h00;
assign TX_DATA_41_const_net_27             = 8'h00;
assign TX_DATA_42_const_net_27             = 8'h00;
assign TX_DATA_43_const_net_27             = 8'h00;
assign TX_DATA_44_const_net_27             = 8'h00;
assign TX_DATA_45_const_net_27             = 8'h00;
assign TX_DATA_46_const_net_27             = 8'h00;
assign TX_DATA_47_const_net_27             = 8'h00;
assign TX_DATA_48_const_net_27             = 8'h00;
assign TX_DATA_49_const_net_27             = 8'h00;
assign TX_DATA_50_const_net_27             = 8'h00;
assign TX_DATA_51_const_net_27             = 8'h00;
assign TX_DATA_52_const_net_27             = 8'h00;
assign TX_DATA_53_const_net_27             = 8'h00;
assign TX_DATA_54_const_net_27             = 8'h00;
assign TX_DATA_55_const_net_27             = 8'h00;
assign TX_DATA_56_const_net_27             = 8'h00;
assign TX_DATA_57_const_net_27             = 8'h00;
assign TX_DATA_58_const_net_27             = 8'h00;
assign TX_DATA_59_const_net_27             = 8'h00;
assign TX_DATA_60_const_net_27             = 8'h00;
assign TX_DATA_61_const_net_27             = 8'h00;
assign TX_DATA_62_const_net_27             = 8'h00;
assign TX_DATA_63_const_net_27             = 8'h00;
assign TX_DATA_64_const_net_27             = 8'h00;
assign TX_DATA_65_const_net_27             = 8'h00;
assign TX_DATA_66_const_net_27             = 8'h00;
assign TX_DATA_67_const_net_27             = 8'h00;
assign TX_DATA_68_const_net_27             = 8'h00;
assign TX_DATA_69_const_net_27             = 8'h00;
assign TX_DATA_70_const_net_27             = 8'h00;
assign TX_DATA_71_const_net_27             = 8'h00;
assign TX_DATA_72_const_net_27             = 8'h00;
assign TX_DATA_73_const_net_27             = 8'h00;
assign TX_DATA_74_const_net_27             = 8'h00;
assign TX_DATA_75_const_net_27             = 8'h00;
assign TX_DATA_76_const_net_27             = 8'h00;
assign TX_DATA_77_const_net_27             = 8'h00;
assign TX_DATA_78_const_net_27             = 8'h00;
assign TX_DATA_79_const_net_27             = 8'h00;
assign TX_DATA_80_const_net_27             = 8'h00;
assign TX_DATA_81_const_net_27             = 8'h00;
assign TX_DATA_82_const_net_27             = 8'h00;
assign TX_DATA_83_const_net_27             = 8'h00;
assign TX_DATA_84_const_net_27             = 8'h00;
assign TX_DATA_85_const_net_27             = 8'h00;
assign TX_DATA_86_const_net_27             = 8'h00;
assign TX_DATA_87_const_net_27             = 8'h00;
assign TX_DATA_88_const_net_27             = 8'h00;
assign TX_DATA_89_const_net_27             = 8'h00;
assign TX_DATA_90_const_net_27             = 8'h00;
assign TX_DATA_91_const_net_27             = 8'h00;
assign TX_DATA_92_const_net_27             = 8'h00;
assign TX_DATA_93_const_net_27             = 8'h00;
assign TX_DATA_94_const_net_27             = 8'h00;
assign TX_DATA_95_const_net_27             = 8'h00;
assign TX_DATA_96_const_net_27             = 8'h00;
assign TX_DATA_97_const_net_27             = 8'h00;
assign TX_DATA_98_const_net_27             = 8'h00;
assign TX_DATA_99_const_net_27             = 8'h00;
assign TX_DATA_100_const_net_27            = 8'h00;
assign TX_DATA_101_const_net_27            = 8'h00;
assign TX_DATA_102_const_net_27            = 8'h00;
assign TX_DATA_103_const_net_27            = 8'h00;
assign TX_DATA_104_const_net_27            = 8'h00;
assign TX_DATA_105_const_net_27            = 8'h00;
assign TX_DATA_106_const_net_27            = 8'h00;
assign TX_DATA_107_const_net_27            = 8'h00;
assign TX_DATA_108_const_net_27            = 8'h00;
assign TX_DATA_109_const_net_27            = 8'h00;
assign TX_DATA_110_const_net_27            = 8'h00;
assign TX_DATA_111_const_net_27            = 8'h00;
assign TX_DATA_112_const_net_27            = 8'h00;
assign TX_DATA_113_const_net_27            = 8'h00;
assign TX_DATA_114_const_net_27            = 8'h00;
assign TX_DATA_115_const_net_27            = 8'h00;
assign TX_DATA_116_const_net_27            = 8'h00;
assign TX_DATA_117_const_net_27            = 8'h00;
assign TX_DATA_118_const_net_27            = 8'h00;
assign TX_DATA_119_const_net_27            = 8'h00;
assign TX_DATA_120_const_net_27            = 8'h00;
assign TX_DATA_121_const_net_27            = 8'h00;
assign TX_DATA_122_const_net_27            = 8'h00;
assign TX_DATA_123_const_net_27            = 8'h00;
assign TX_DATA_124_const_net_27            = 8'h00;
assign TX_DATA_125_const_net_27            = 8'h00;
assign TX_DATA_126_const_net_27            = 8'h00;
assign TX_DATA_127_const_net_27            = 8'h00;
assign OE_DATA_1_const_net_24              = 4'h0;
assign OE_DATA_2_const_net_24              = 4'h0;
assign OE_DATA_3_const_net_24              = 4'h0;
assign OE_DATA_4_const_net_24              = 4'h0;
assign OE_DATA_5_const_net_24              = 4'h0;
assign OE_DATA_6_const_net_24              = 4'h0;
assign OE_DATA_7_const_net_24              = 4'h0;
assign OE_DATA_8_const_net_27              = 4'h0;
assign OE_DATA_9_const_net_27              = 4'h0;
assign OE_DATA_10_const_net_27             = 4'h0;
assign OE_DATA_11_const_net_27             = 4'h0;
assign OE_DATA_12_const_net_27             = 4'h0;
assign OE_DATA_13_const_net_27             = 4'h0;
assign OE_DATA_14_const_net_27             = 4'h0;
assign OE_DATA_15_const_net_27             = 4'h0;
assign OE_DATA_16_const_net_27             = 4'h0;
assign OE_DATA_17_const_net_27             = 4'h0;
assign OE_DATA_18_const_net_27             = 4'h0;
assign OE_DATA_19_const_net_27             = 4'h0;
assign OE_DATA_20_const_net_27             = 4'h0;
assign OE_DATA_21_const_net_27             = 4'h0;
assign OE_DATA_22_const_net_27             = 4'h0;
assign OE_DATA_23_const_net_27             = 4'h0;
assign OE_DATA_24_const_net_27             = 4'h0;
assign OE_DATA_25_const_net_27             = 4'h0;
assign OE_DATA_26_const_net_27             = 4'h0;
assign OE_DATA_27_const_net_27             = 4'h0;
assign OE_DATA_28_const_net_27             = 4'h0;
assign OE_DATA_29_const_net_27             = 4'h0;
assign OE_DATA_30_const_net_27             = 4'h0;
assign OE_DATA_31_const_net_27             = 4'h0;
assign OE_DATA_32_const_net_27             = 4'h0;
assign OE_DATA_33_const_net_27             = 4'h0;
assign OE_DATA_34_const_net_27             = 4'h0;
assign OE_DATA_35_const_net_27             = 4'h0;
assign OE_DATA_36_const_net_27             = 4'h0;
assign OE_DATA_37_const_net_27             = 4'h0;
assign OE_DATA_38_const_net_27             = 4'h0;
assign OE_DATA_39_const_net_27             = 4'h0;
assign OE_DATA_40_const_net_27             = 4'h0;
assign OE_DATA_41_const_net_27             = 4'h0;
assign OE_DATA_42_const_net_27             = 4'h0;
assign OE_DATA_43_const_net_27             = 4'h0;
assign OE_DATA_44_const_net_27             = 4'h0;
assign OE_DATA_45_const_net_27             = 4'h0;
assign OE_DATA_46_const_net_27             = 4'h0;
assign OE_DATA_47_const_net_27             = 4'h0;
assign OE_DATA_48_const_net_27             = 4'h0;
assign OE_DATA_49_const_net_27             = 4'h0;
assign OE_DATA_50_const_net_27             = 4'h0;
assign OE_DATA_51_const_net_27             = 4'h0;
assign OE_DATA_52_const_net_27             = 4'h0;
assign OE_DATA_53_const_net_27             = 4'h0;
assign OE_DATA_54_const_net_27             = 4'h0;
assign OE_DATA_55_const_net_27             = 4'h0;
assign OE_DATA_56_const_net_27             = 4'h0;
assign OE_DATA_57_const_net_27             = 4'h0;
assign OE_DATA_58_const_net_27             = 4'h0;
assign OE_DATA_59_const_net_27             = 4'h0;
assign OE_DATA_60_const_net_27             = 4'h0;
assign OE_DATA_61_const_net_27             = 4'h0;
assign OE_DATA_62_const_net_27             = 4'h0;
assign OE_DATA_63_const_net_27             = 4'h0;
assign OE_DATA_64_const_net_27             = 4'h0;
assign OE_DATA_65_const_net_27             = 4'h0;
assign OE_DATA_66_const_net_27             = 4'h0;
assign OE_DATA_67_const_net_27             = 4'h0;
assign OE_DATA_68_const_net_27             = 4'h0;
assign OE_DATA_69_const_net_27             = 4'h0;
assign OE_DATA_70_const_net_27             = 4'h0;
assign OE_DATA_71_const_net_27             = 4'h0;
assign OE_DATA_72_const_net_27             = 4'h0;
assign OE_DATA_73_const_net_27             = 4'h0;
assign OE_DATA_74_const_net_27             = 4'h0;
assign OE_DATA_75_const_net_27             = 4'h0;
assign OE_DATA_76_const_net_27             = 4'h0;
assign OE_DATA_77_const_net_27             = 4'h0;
assign OE_DATA_78_const_net_27             = 4'h0;
assign OE_DATA_79_const_net_27             = 4'h0;
assign OE_DATA_80_const_net_27             = 4'h0;
assign OE_DATA_81_const_net_27             = 4'h0;
assign OE_DATA_82_const_net_27             = 4'h0;
assign OE_DATA_83_const_net_27             = 4'h0;
assign OE_DATA_84_const_net_27             = 4'h0;
assign OE_DATA_85_const_net_27             = 4'h0;
assign OE_DATA_86_const_net_27             = 4'h0;
assign OE_DATA_87_const_net_27             = 4'h0;
assign OE_DATA_88_const_net_27             = 4'h0;
assign OE_DATA_89_const_net_27             = 4'h0;
assign OE_DATA_90_const_net_27             = 4'h0;
assign OE_DATA_91_const_net_27             = 4'h0;
assign OE_DATA_92_const_net_27             = 4'h0;
assign OE_DATA_93_const_net_27             = 4'h0;
assign OE_DATA_94_const_net_27             = 4'h0;
assign OE_DATA_95_const_net_27             = 4'h0;
assign OE_DATA_96_const_net_27             = 4'h0;
assign OE_DATA_97_const_net_27             = 4'h0;
assign OE_DATA_98_const_net_27             = 4'h0;
assign OE_DATA_99_const_net_27             = 4'h0;
assign OE_DATA_100_const_net_27            = 4'h0;
assign OE_DATA_101_const_net_27            = 4'h0;
assign OE_DATA_102_const_net_27            = 4'h0;
assign OE_DATA_103_const_net_27            = 4'h0;
assign OE_DATA_104_const_net_27            = 4'h0;
assign OE_DATA_105_const_net_27            = 4'h0;
assign OE_DATA_106_const_net_27            = 4'h0;
assign OE_DATA_107_const_net_27            = 4'h0;
assign OE_DATA_108_const_net_27            = 4'h0;
assign OE_DATA_109_const_net_27            = 4'h0;
assign OE_DATA_110_const_net_27            = 4'h0;
assign OE_DATA_111_const_net_27            = 4'h0;
assign OE_DATA_112_const_net_27            = 4'h0;
assign OE_DATA_113_const_net_27            = 4'h0;
assign OE_DATA_114_const_net_27            = 4'h0;
assign OE_DATA_115_const_net_27            = 4'h0;
assign OE_DATA_116_const_net_27            = 4'h0;
assign OE_DATA_117_const_net_27            = 4'h0;
assign OE_DATA_118_const_net_27            = 4'h0;
assign OE_DATA_119_const_net_27            = 4'h0;
assign OE_DATA_120_const_net_27            = 4'h0;
assign OE_DATA_121_const_net_27            = 4'h0;
assign OE_DATA_122_const_net_27            = 4'h0;
assign OE_DATA_123_const_net_27            = 4'h0;
assign OE_DATA_124_const_net_27            = 4'h0;
assign OE_DATA_125_const_net_27            = 4'h0;
assign OE_DATA_126_const_net_27            = 4'h0;
assign OE_DATA_127_const_net_27            = 4'h0;
assign RX_DQS_90_const_net_19              = 2'h0;
assign FIFO_WR_PTR_const_net_20            = 3'h0;
assign FIFO_RD_PTR_const_net_20            = 3'h0;
assign EYE_MONITOR_LANE_WIDTH_const_net_22 = 3'h0;
assign TX_DATA_1_const_net_22              = 2'h0;
assign TX_DATA_2_const_net_24              = 2'h0;
assign TX_DATA_3_const_net_24              = 2'h0;
assign TX_DATA_4_const_net_24              = 2'h0;
assign TX_DATA_5_const_net_24              = 2'h0;
assign TX_DATA_6_const_net_24              = 2'h0;
assign TX_DATA_7_const_net_24              = 2'h0;
assign TX_DATA_8_const_net_27              = 2'h0;
assign TX_DATA_9_const_net_27              = 2'h0;
assign TX_DATA_10_const_net_27             = 2'h0;
assign TX_DATA_11_const_net_27             = 2'h0;
assign TX_DATA_12_const_net_28             = 2'h0;
assign TX_DATA_13_const_net_28             = 2'h0;
assign TX_DATA_14_const_net_28             = 2'h0;
assign TX_DATA_15_const_net_28             = 2'h0;
assign TX_DATA_16_const_net_28             = 2'h0;
assign TX_DATA_17_const_net_28             = 2'h0;
assign TX_DATA_18_const_net_28             = 2'h0;
assign TX_DATA_19_const_net_28             = 2'h0;
assign TX_DATA_20_const_net_28             = 2'h0;
assign TX_DATA_21_const_net_28             = 2'h0;
assign TX_DATA_22_const_net_28             = 2'h0;
assign TX_DATA_23_const_net_28             = 2'h0;
assign TX_DATA_24_const_net_28             = 2'h0;
assign TX_DATA_25_const_net_28             = 2'h0;
assign TX_DATA_26_const_net_28             = 2'h0;
assign TX_DATA_27_const_net_28             = 2'h0;
assign TX_DATA_28_const_net_28             = 2'h0;
assign TX_DATA_29_const_net_28             = 2'h0;
assign TX_DATA_30_const_net_28             = 2'h0;
assign TX_DATA_31_const_net_28             = 2'h0;
assign TX_DATA_32_const_net_28             = 2'h0;
assign TX_DATA_33_const_net_28             = 2'h0;
assign TX_DATA_34_const_net_28             = 2'h0;
assign TX_DATA_35_const_net_28             = 2'h0;
assign TX_DATA_36_const_net_28             = 2'h0;
assign TX_DATA_37_const_net_28             = 2'h0;
assign TX_DATA_38_const_net_28             = 2'h0;
assign TX_DATA_39_const_net_28             = 2'h0;
assign TX_DATA_40_const_net_28             = 2'h0;
assign TX_DATA_41_const_net_28             = 2'h0;
assign TX_DATA_42_const_net_28             = 2'h0;
assign TX_DATA_43_const_net_28             = 2'h0;
assign TX_DATA_44_const_net_28             = 2'h0;
assign TX_DATA_45_const_net_28             = 2'h0;
assign TX_DATA_46_const_net_28             = 2'h0;
assign TX_DATA_47_const_net_28             = 2'h0;
assign TX_DATA_48_const_net_28             = 2'h0;
assign TX_DATA_49_const_net_28             = 2'h0;
assign TX_DATA_50_const_net_28             = 2'h0;
assign TX_DATA_51_const_net_28             = 2'h0;
assign TX_DATA_52_const_net_28             = 2'h0;
assign TX_DATA_53_const_net_28             = 2'h0;
assign TX_DATA_54_const_net_28             = 2'h0;
assign TX_DATA_55_const_net_28             = 2'h0;
assign TX_DATA_56_const_net_28             = 2'h0;
assign TX_DATA_57_const_net_28             = 2'h0;
assign TX_DATA_58_const_net_28             = 2'h0;
assign TX_DATA_59_const_net_28             = 2'h0;
assign TX_DATA_60_const_net_28             = 2'h0;
assign TX_DATA_61_const_net_28             = 2'h0;
assign TX_DATA_62_const_net_28             = 2'h0;
assign TX_DATA_63_const_net_28             = 2'h0;
assign TX_DATA_64_const_net_28             = 2'h0;
assign TX_DATA_65_const_net_28             = 2'h0;
assign TX_DATA_66_const_net_28             = 2'h0;
assign TX_DATA_67_const_net_28             = 2'h0;
assign TX_DATA_68_const_net_28             = 2'h0;
assign TX_DATA_69_const_net_28             = 2'h0;
assign TX_DATA_70_const_net_28             = 2'h0;
assign TX_DATA_71_const_net_28             = 2'h0;
assign TX_DATA_72_const_net_28             = 2'h0;
assign TX_DATA_73_const_net_28             = 2'h0;
assign TX_DATA_74_const_net_28             = 2'h0;
assign TX_DATA_75_const_net_28             = 2'h0;
assign TX_DATA_76_const_net_28             = 2'h0;
assign TX_DATA_77_const_net_28             = 2'h0;
assign TX_DATA_78_const_net_28             = 2'h0;
assign TX_DATA_79_const_net_28             = 2'h0;
assign TX_DATA_80_const_net_28             = 2'h0;
assign TX_DATA_81_const_net_28             = 2'h0;
assign TX_DATA_82_const_net_28             = 2'h0;
assign TX_DATA_83_const_net_28             = 2'h0;
assign TX_DATA_84_const_net_28             = 2'h0;
assign TX_DATA_85_const_net_28             = 2'h0;
assign TX_DATA_86_const_net_28             = 2'h0;
assign TX_DATA_87_const_net_28             = 2'h0;
assign TX_DATA_88_const_net_28             = 2'h0;
assign TX_DATA_89_const_net_28             = 2'h0;
assign TX_DATA_90_const_net_28             = 2'h0;
assign TX_DATA_91_const_net_28             = 2'h0;
assign TX_DATA_92_const_net_28             = 2'h0;
assign TX_DATA_93_const_net_28             = 2'h0;
assign TX_DATA_94_const_net_28             = 2'h0;
assign TX_DATA_95_const_net_28             = 2'h0;
assign TX_DATA_96_const_net_28             = 2'h0;
assign TX_DATA_97_const_net_28             = 2'h0;
assign TX_DATA_98_const_net_28             = 2'h0;
assign TX_DATA_99_const_net_28             = 2'h0;
assign TX_DATA_100_const_net_28            = 2'h0;
assign TX_DATA_101_const_net_28            = 2'h0;
assign TX_DATA_102_const_net_28            = 2'h0;
assign TX_DATA_103_const_net_28            = 2'h0;
assign TX_DATA_104_const_net_28            = 2'h0;
assign TX_DATA_105_const_net_28            = 2'h0;
assign TX_DATA_106_const_net_28            = 2'h0;
assign TX_DATA_107_const_net_28            = 2'h0;
assign TX_DATA_108_const_net_28            = 2'h0;
assign TX_DATA_109_const_net_28            = 2'h0;
assign TX_DATA_110_const_net_28            = 2'h0;
assign TX_DATA_111_const_net_28            = 2'h0;
assign TX_DATA_112_const_net_28            = 2'h0;
assign TX_DATA_113_const_net_28            = 2'h0;
assign TX_DATA_114_const_net_28            = 2'h0;
assign TX_DATA_115_const_net_28            = 2'h0;
assign TX_DATA_116_const_net_28            = 2'h0;
assign TX_DATA_117_const_net_28            = 2'h0;
assign TX_DATA_118_const_net_28            = 2'h0;
assign TX_DATA_119_const_net_28            = 2'h0;
assign TX_DATA_120_const_net_28            = 2'h0;
assign TX_DATA_121_const_net_28            = 2'h0;
assign TX_DATA_122_const_net_28            = 2'h0;
assign TX_DATA_123_const_net_28            = 2'h0;
assign TX_DATA_124_const_net_28            = 2'h0;
assign TX_DATA_125_const_net_28            = 2'h0;
assign TX_DATA_126_const_net_28            = 2'h0;
assign TX_DATA_127_const_net_28            = 2'h0;
assign OE_DATA_1_const_net_25              = 2'h0;
assign OE_DATA_2_const_net_25              = 2'h0;
assign OE_DATA_3_const_net_25              = 2'h0;
assign OE_DATA_4_const_net_25              = 2'h0;
assign OE_DATA_5_const_net_25              = 2'h0;
assign OE_DATA_6_const_net_25              = 2'h0;
assign OE_DATA_7_const_net_25              = 2'h0;
assign OE_DATA_8_const_net_28              = 2'h0;
assign OE_DATA_9_const_net_28              = 2'h0;
assign OE_DATA_10_const_net_28             = 2'h0;
assign OE_DATA_11_const_net_28             = 2'h0;
assign OE_DATA_12_const_net_28             = 2'h0;
assign OE_DATA_13_const_net_28             = 2'h0;
assign OE_DATA_14_const_net_28             = 2'h0;
assign OE_DATA_15_const_net_28             = 2'h0;
assign OE_DATA_16_const_net_28             = 2'h0;
assign OE_DATA_17_const_net_28             = 2'h0;
assign OE_DATA_18_const_net_28             = 2'h0;
assign OE_DATA_19_const_net_28             = 2'h0;
assign OE_DATA_20_const_net_28             = 2'h0;
assign OE_DATA_21_const_net_28             = 2'h0;
assign OE_DATA_22_const_net_28             = 2'h0;
assign OE_DATA_23_const_net_28             = 2'h0;
assign OE_DATA_24_const_net_28             = 2'h0;
assign OE_DATA_25_const_net_28             = 2'h0;
assign OE_DATA_26_const_net_28             = 2'h0;
assign OE_DATA_27_const_net_28             = 2'h0;
assign OE_DATA_28_const_net_28             = 2'h0;
assign OE_DATA_29_const_net_28             = 2'h0;
assign OE_DATA_30_const_net_28             = 2'h0;
assign OE_DATA_31_const_net_28             = 2'h0;
assign OE_DATA_32_const_net_28             = 2'h0;
assign OE_DATA_33_const_net_28             = 2'h0;
assign OE_DATA_34_const_net_28             = 2'h0;
assign OE_DATA_35_const_net_28             = 2'h0;
assign OE_DATA_36_const_net_28             = 2'h0;
assign OE_DATA_37_const_net_28             = 2'h0;
assign OE_DATA_38_const_net_28             = 2'h0;
assign OE_DATA_39_const_net_28             = 2'h0;
assign OE_DATA_40_const_net_28             = 2'h0;
assign OE_DATA_41_const_net_28             = 2'h0;
assign OE_DATA_42_const_net_28             = 2'h0;
assign OE_DATA_43_const_net_28             = 2'h0;
assign OE_DATA_44_const_net_28             = 2'h0;
assign OE_DATA_45_const_net_28             = 2'h0;
assign OE_DATA_46_const_net_28             = 2'h0;
assign OE_DATA_47_const_net_28             = 2'h0;
assign OE_DATA_48_const_net_28             = 2'h0;
assign OE_DATA_49_const_net_28             = 2'h0;
assign OE_DATA_50_const_net_28             = 2'h0;
assign OE_DATA_51_const_net_28             = 2'h0;
assign OE_DATA_52_const_net_28             = 2'h0;
assign OE_DATA_53_const_net_28             = 2'h0;
assign OE_DATA_54_const_net_28             = 2'h0;
assign OE_DATA_55_const_net_28             = 2'h0;
assign OE_DATA_56_const_net_28             = 2'h0;
assign OE_DATA_57_const_net_28             = 2'h0;
assign OE_DATA_58_const_net_28             = 2'h0;
assign OE_DATA_59_const_net_28             = 2'h0;
assign OE_DATA_60_const_net_28             = 2'h0;
assign OE_DATA_61_const_net_28             = 2'h0;
assign OE_DATA_62_const_net_28             = 2'h0;
assign OE_DATA_63_const_net_28             = 2'h0;
assign OE_DATA_64_const_net_28             = 2'h0;
assign OE_DATA_65_const_net_28             = 2'h0;
assign OE_DATA_66_const_net_28             = 2'h0;
assign OE_DATA_67_const_net_28             = 2'h0;
assign OE_DATA_68_const_net_28             = 2'h0;
assign OE_DATA_69_const_net_28             = 2'h0;
assign OE_DATA_70_const_net_28             = 2'h0;
assign OE_DATA_71_const_net_28             = 2'h0;
assign OE_DATA_72_const_net_28             = 2'h0;
assign OE_DATA_73_const_net_28             = 2'h0;
assign OE_DATA_74_const_net_28             = 2'h0;
assign OE_DATA_75_const_net_28             = 2'h0;
assign OE_DATA_76_const_net_28             = 2'h0;
assign OE_DATA_77_const_net_28             = 2'h0;
assign OE_DATA_78_const_net_28             = 2'h0;
assign OE_DATA_79_const_net_28             = 2'h0;
assign OE_DATA_80_const_net_28             = 2'h0;
assign OE_DATA_81_const_net_28             = 2'h0;
assign OE_DATA_82_const_net_28             = 2'h0;
assign OE_DATA_83_const_net_28             = 2'h0;
assign OE_DATA_84_const_net_28             = 2'h0;
assign OE_DATA_85_const_net_28             = 2'h0;
assign OE_DATA_86_const_net_28             = 2'h0;
assign OE_DATA_87_const_net_28             = 2'h0;
assign OE_DATA_88_const_net_28             = 2'h0;
assign OE_DATA_89_const_net_28             = 2'h0;
assign OE_DATA_90_const_net_28             = 2'h0;
assign OE_DATA_91_const_net_28             = 2'h0;
assign OE_DATA_92_const_net_28             = 2'h0;
assign OE_DATA_93_const_net_28             = 2'h0;
assign OE_DATA_94_const_net_28             = 2'h0;
assign OE_DATA_95_const_net_28             = 2'h0;
assign OE_DATA_96_const_net_28             = 2'h0;
assign OE_DATA_97_const_net_28             = 2'h0;
assign OE_DATA_98_const_net_28             = 2'h0;
assign OE_DATA_99_const_net_28             = 2'h0;
assign OE_DATA_100_const_net_28            = 2'h0;
assign OE_DATA_101_const_net_28            = 2'h0;
assign OE_DATA_102_const_net_28            = 2'h0;
assign OE_DATA_103_const_net_28            = 2'h0;
assign OE_DATA_104_const_net_28            = 2'h0;
assign OE_DATA_105_const_net_28            = 2'h0;
assign OE_DATA_106_const_net_28            = 2'h0;
assign OE_DATA_107_const_net_28            = 2'h0;
assign OE_DATA_108_const_net_28            = 2'h0;
assign OE_DATA_109_const_net_28            = 2'h0;
assign OE_DATA_110_const_net_28            = 2'h0;
assign OE_DATA_111_const_net_28            = 2'h0;
assign OE_DATA_112_const_net_28            = 2'h0;
assign OE_DATA_113_const_net_28            = 2'h0;
assign OE_DATA_114_const_net_28            = 2'h0;
assign OE_DATA_115_const_net_28            = 2'h0;
assign OE_DATA_116_const_net_28            = 2'h0;
assign OE_DATA_117_const_net_28            = 2'h0;
assign OE_DATA_118_const_net_28            = 2'h0;
assign OE_DATA_119_const_net_28            = 2'h0;
assign OE_DATA_120_const_net_28            = 2'h0;
assign OE_DATA_121_const_net_28            = 2'h0;
assign OE_DATA_122_const_net_28            = 2'h0;
assign OE_DATA_123_const_net_28            = 2'h0;
assign OE_DATA_124_const_net_28            = 2'h0;
assign OE_DATA_125_const_net_28            = 2'h0;
assign OE_DATA_126_const_net_28            = 2'h0;
assign OE_DATA_127_const_net_28            = 2'h0;
assign RX_DQS_90_const_net_20              = 2'h0;
assign EYE_MONITOR_LANE_WIDTH_const_net_23 = 3'h0;
assign TX_DATA_1_const_net_23              = 8'h00;
assign TX_DATA_2_const_net_25              = 8'h00;
assign TX_DATA_3_const_net_25              = 8'h00;
assign TX_DATA_4_const_net_25              = 8'h00;
assign TX_DATA_5_const_net_25              = 8'h00;
assign TX_DATA_6_const_net_25              = 8'h00;
assign TX_DATA_7_const_net_25              = 8'h00;
assign TX_DATA_8_const_net_28              = 8'h00;
assign TX_DATA_9_const_net_28              = 8'h00;
assign TX_DATA_10_const_net_28             = 8'h00;
assign TX_DATA_11_const_net_28             = 8'h00;
assign TX_DATA_12_const_net_29             = 8'h00;
assign TX_DATA_13_const_net_29             = 8'h00;
assign TX_DATA_14_const_net_29             = 8'h00;
assign TX_DATA_15_const_net_29             = 8'h00;
assign TX_DATA_16_const_net_29             = 8'h00;
assign TX_DATA_17_const_net_29             = 8'h00;
assign TX_DATA_18_const_net_29             = 8'h00;
assign TX_DATA_19_const_net_29             = 8'h00;
assign TX_DATA_20_const_net_29             = 8'h00;
assign TX_DATA_21_const_net_29             = 8'h00;
assign TX_DATA_22_const_net_29             = 8'h00;
assign TX_DATA_23_const_net_29             = 8'h00;
assign TX_DATA_24_const_net_29             = 8'h00;
assign TX_DATA_25_const_net_29             = 8'h00;
assign TX_DATA_26_const_net_29             = 8'h00;
assign TX_DATA_27_const_net_29             = 8'h00;
assign TX_DATA_28_const_net_29             = 8'h00;
assign TX_DATA_29_const_net_29             = 8'h00;
assign TX_DATA_30_const_net_29             = 8'h00;
assign TX_DATA_31_const_net_29             = 8'h00;
assign TX_DATA_32_const_net_29             = 8'h00;
assign TX_DATA_33_const_net_29             = 8'h00;
assign TX_DATA_34_const_net_29             = 8'h00;
assign TX_DATA_35_const_net_29             = 8'h00;
assign TX_DATA_36_const_net_29             = 8'h00;
assign TX_DATA_37_const_net_29             = 8'h00;
assign TX_DATA_38_const_net_29             = 8'h00;
assign TX_DATA_39_const_net_29             = 8'h00;
assign TX_DATA_40_const_net_29             = 8'h00;
assign TX_DATA_41_const_net_29             = 8'h00;
assign TX_DATA_42_const_net_29             = 8'h00;
assign TX_DATA_43_const_net_29             = 8'h00;
assign TX_DATA_44_const_net_29             = 8'h00;
assign TX_DATA_45_const_net_29             = 8'h00;
assign TX_DATA_46_const_net_29             = 8'h00;
assign TX_DATA_47_const_net_29             = 8'h00;
assign TX_DATA_48_const_net_29             = 8'h00;
assign TX_DATA_49_const_net_29             = 8'h00;
assign TX_DATA_50_const_net_29             = 8'h00;
assign TX_DATA_51_const_net_29             = 8'h00;
assign TX_DATA_52_const_net_29             = 8'h00;
assign TX_DATA_53_const_net_29             = 8'h00;
assign TX_DATA_54_const_net_29             = 8'h00;
assign TX_DATA_55_const_net_29             = 8'h00;
assign TX_DATA_56_const_net_29             = 8'h00;
assign TX_DATA_57_const_net_29             = 8'h00;
assign TX_DATA_58_const_net_29             = 8'h00;
assign TX_DATA_59_const_net_29             = 8'h00;
assign TX_DATA_60_const_net_29             = 8'h00;
assign TX_DATA_61_const_net_29             = 8'h00;
assign TX_DATA_62_const_net_29             = 8'h00;
assign TX_DATA_63_const_net_29             = 8'h00;
assign TX_DATA_64_const_net_29             = 8'h00;
assign TX_DATA_65_const_net_29             = 8'h00;
assign TX_DATA_66_const_net_29             = 8'h00;
assign TX_DATA_67_const_net_29             = 8'h00;
assign TX_DATA_68_const_net_29             = 8'h00;
assign TX_DATA_69_const_net_29             = 8'h00;
assign TX_DATA_70_const_net_29             = 8'h00;
assign TX_DATA_71_const_net_29             = 8'h00;
assign TX_DATA_72_const_net_29             = 8'h00;
assign TX_DATA_73_const_net_29             = 8'h00;
assign TX_DATA_74_const_net_29             = 8'h00;
assign TX_DATA_75_const_net_29             = 8'h00;
assign TX_DATA_76_const_net_29             = 8'h00;
assign TX_DATA_77_const_net_29             = 8'h00;
assign TX_DATA_78_const_net_29             = 8'h00;
assign TX_DATA_79_const_net_29             = 8'h00;
assign TX_DATA_80_const_net_29             = 8'h00;
assign TX_DATA_81_const_net_29             = 8'h00;
assign TX_DATA_82_const_net_29             = 8'h00;
assign TX_DATA_83_const_net_29             = 8'h00;
assign TX_DATA_84_const_net_29             = 8'h00;
assign TX_DATA_85_const_net_29             = 8'h00;
assign TX_DATA_86_const_net_29             = 8'h00;
assign TX_DATA_87_const_net_29             = 8'h00;
assign TX_DATA_88_const_net_29             = 8'h00;
assign TX_DATA_89_const_net_29             = 8'h00;
assign TX_DATA_90_const_net_29             = 8'h00;
assign TX_DATA_91_const_net_29             = 8'h00;
assign TX_DATA_92_const_net_29             = 8'h00;
assign TX_DATA_93_const_net_29             = 8'h00;
assign TX_DATA_94_const_net_29             = 8'h00;
assign TX_DATA_95_const_net_29             = 8'h00;
assign TX_DATA_96_const_net_29             = 8'h00;
assign TX_DATA_97_const_net_29             = 8'h00;
assign TX_DATA_98_const_net_29             = 8'h00;
assign TX_DATA_99_const_net_29             = 8'h00;
assign TX_DATA_100_const_net_29            = 8'h00;
assign TX_DATA_101_const_net_29            = 8'h00;
assign TX_DATA_102_const_net_29            = 8'h00;
assign TX_DATA_103_const_net_29            = 8'h00;
assign TX_DATA_104_const_net_29            = 8'h00;
assign TX_DATA_105_const_net_29            = 8'h00;
assign TX_DATA_106_const_net_29            = 8'h00;
assign TX_DATA_107_const_net_29            = 8'h00;
assign TX_DATA_108_const_net_29            = 8'h00;
assign TX_DATA_109_const_net_29            = 8'h00;
assign TX_DATA_110_const_net_29            = 8'h00;
assign TX_DATA_111_const_net_29            = 8'h00;
assign TX_DATA_112_const_net_29            = 8'h00;
assign TX_DATA_113_const_net_29            = 8'h00;
assign TX_DATA_114_const_net_29            = 8'h00;
assign TX_DATA_115_const_net_29            = 8'h00;
assign TX_DATA_116_const_net_29            = 8'h00;
assign TX_DATA_117_const_net_29            = 8'h00;
assign TX_DATA_118_const_net_29            = 8'h00;
assign TX_DATA_119_const_net_29            = 8'h00;
assign TX_DATA_120_const_net_29            = 8'h00;
assign TX_DATA_121_const_net_29            = 8'h00;
assign TX_DATA_122_const_net_29            = 8'h00;
assign TX_DATA_123_const_net_29            = 8'h00;
assign TX_DATA_124_const_net_29            = 8'h00;
assign TX_DATA_125_const_net_29            = 8'h00;
assign TX_DATA_126_const_net_29            = 8'h00;
assign TX_DATA_127_const_net_29            = 8'h00;
assign OE_DATA_1_const_net_26              = 4'h0;
assign OE_DATA_2_const_net_26              = 4'h0;
assign OE_DATA_3_const_net_26              = 4'h0;
assign OE_DATA_4_const_net_26              = 4'h0;
assign OE_DATA_5_const_net_26              = 4'h0;
assign OE_DATA_6_const_net_26              = 4'h0;
assign OE_DATA_7_const_net_26              = 4'h0;
assign OE_DATA_8_const_net_29              = 4'h0;
assign OE_DATA_9_const_net_29              = 4'h0;
assign OE_DATA_10_const_net_29             = 4'h0;
assign OE_DATA_11_const_net_29             = 4'h0;
assign OE_DATA_12_const_net_29             = 4'h0;
assign OE_DATA_13_const_net_29             = 4'h0;
assign OE_DATA_14_const_net_29             = 4'h0;
assign OE_DATA_15_const_net_29             = 4'h0;
assign OE_DATA_16_const_net_29             = 4'h0;
assign OE_DATA_17_const_net_29             = 4'h0;
assign OE_DATA_18_const_net_29             = 4'h0;
assign OE_DATA_19_const_net_29             = 4'h0;
assign OE_DATA_20_const_net_29             = 4'h0;
assign OE_DATA_21_const_net_29             = 4'h0;
assign OE_DATA_22_const_net_29             = 4'h0;
assign OE_DATA_23_const_net_29             = 4'h0;
assign OE_DATA_24_const_net_29             = 4'h0;
assign OE_DATA_25_const_net_29             = 4'h0;
assign OE_DATA_26_const_net_29             = 4'h0;
assign OE_DATA_27_const_net_29             = 4'h0;
assign OE_DATA_28_const_net_29             = 4'h0;
assign OE_DATA_29_const_net_29             = 4'h0;
assign OE_DATA_30_const_net_29             = 4'h0;
assign OE_DATA_31_const_net_29             = 4'h0;
assign OE_DATA_32_const_net_29             = 4'h0;
assign OE_DATA_33_const_net_29             = 4'h0;
assign OE_DATA_34_const_net_29             = 4'h0;
assign OE_DATA_35_const_net_29             = 4'h0;
assign OE_DATA_36_const_net_29             = 4'h0;
assign OE_DATA_37_const_net_29             = 4'h0;
assign OE_DATA_38_const_net_29             = 4'h0;
assign OE_DATA_39_const_net_29             = 4'h0;
assign OE_DATA_40_const_net_29             = 4'h0;
assign OE_DATA_41_const_net_29             = 4'h0;
assign OE_DATA_42_const_net_29             = 4'h0;
assign OE_DATA_43_const_net_29             = 4'h0;
assign OE_DATA_44_const_net_29             = 4'h0;
assign OE_DATA_45_const_net_29             = 4'h0;
assign OE_DATA_46_const_net_29             = 4'h0;
assign OE_DATA_47_const_net_29             = 4'h0;
assign OE_DATA_48_const_net_29             = 4'h0;
assign OE_DATA_49_const_net_29             = 4'h0;
assign OE_DATA_50_const_net_29             = 4'h0;
assign OE_DATA_51_const_net_29             = 4'h0;
assign OE_DATA_52_const_net_29             = 4'h0;
assign OE_DATA_53_const_net_29             = 4'h0;
assign OE_DATA_54_const_net_29             = 4'h0;
assign OE_DATA_55_const_net_29             = 4'h0;
assign OE_DATA_56_const_net_29             = 4'h0;
assign OE_DATA_57_const_net_29             = 4'h0;
assign OE_DATA_58_const_net_29             = 4'h0;
assign OE_DATA_59_const_net_29             = 4'h0;
assign OE_DATA_60_const_net_29             = 4'h0;
assign OE_DATA_61_const_net_29             = 4'h0;
assign OE_DATA_62_const_net_29             = 4'h0;
assign OE_DATA_63_const_net_29             = 4'h0;
assign OE_DATA_64_const_net_29             = 4'h0;
assign OE_DATA_65_const_net_29             = 4'h0;
assign OE_DATA_66_const_net_29             = 4'h0;
assign OE_DATA_67_const_net_29             = 4'h0;
assign OE_DATA_68_const_net_29             = 4'h0;
assign OE_DATA_69_const_net_29             = 4'h0;
assign OE_DATA_70_const_net_29             = 4'h0;
assign OE_DATA_71_const_net_29             = 4'h0;
assign OE_DATA_72_const_net_29             = 4'h0;
assign OE_DATA_73_const_net_29             = 4'h0;
assign OE_DATA_74_const_net_29             = 4'h0;
assign OE_DATA_75_const_net_29             = 4'h0;
assign OE_DATA_76_const_net_29             = 4'h0;
assign OE_DATA_77_const_net_29             = 4'h0;
assign OE_DATA_78_const_net_29             = 4'h0;
assign OE_DATA_79_const_net_29             = 4'h0;
assign OE_DATA_80_const_net_29             = 4'h0;
assign OE_DATA_81_const_net_29             = 4'h0;
assign OE_DATA_82_const_net_29             = 4'h0;
assign OE_DATA_83_const_net_29             = 4'h0;
assign OE_DATA_84_const_net_29             = 4'h0;
assign OE_DATA_85_const_net_29             = 4'h0;
assign OE_DATA_86_const_net_29             = 4'h0;
assign OE_DATA_87_const_net_29             = 4'h0;
assign OE_DATA_88_const_net_29             = 4'h0;
assign OE_DATA_89_const_net_29             = 4'h0;
assign OE_DATA_90_const_net_29             = 4'h0;
assign OE_DATA_91_const_net_29             = 4'h0;
assign OE_DATA_92_const_net_29             = 4'h0;
assign OE_DATA_93_const_net_29             = 4'h0;
assign OE_DATA_94_const_net_29             = 4'h0;
assign OE_DATA_95_const_net_29             = 4'h0;
assign OE_DATA_96_const_net_29             = 4'h0;
assign OE_DATA_97_const_net_29             = 4'h0;
assign OE_DATA_98_const_net_29             = 4'h0;
assign OE_DATA_99_const_net_29             = 4'h0;
assign OE_DATA_100_const_net_29            = 4'h0;
assign OE_DATA_101_const_net_29            = 4'h0;
assign OE_DATA_102_const_net_29            = 4'h0;
assign OE_DATA_103_const_net_29            = 4'h0;
assign OE_DATA_104_const_net_29            = 4'h0;
assign OE_DATA_105_const_net_29            = 4'h0;
assign OE_DATA_106_const_net_29            = 4'h0;
assign OE_DATA_107_const_net_29            = 4'h0;
assign OE_DATA_108_const_net_29            = 4'h0;
assign OE_DATA_109_const_net_29            = 4'h0;
assign OE_DATA_110_const_net_29            = 4'h0;
assign OE_DATA_111_const_net_29            = 4'h0;
assign OE_DATA_112_const_net_29            = 4'h0;
assign OE_DATA_113_const_net_29            = 4'h0;
assign OE_DATA_114_const_net_29            = 4'h0;
assign OE_DATA_115_const_net_29            = 4'h0;
assign OE_DATA_116_const_net_29            = 4'h0;
assign OE_DATA_117_const_net_29            = 4'h0;
assign OE_DATA_118_const_net_29            = 4'h0;
assign OE_DATA_119_const_net_29            = 4'h0;
assign OE_DATA_120_const_net_29            = 4'h0;
assign OE_DATA_121_const_net_29            = 4'h0;
assign OE_DATA_122_const_net_29            = 4'h0;
assign OE_DATA_123_const_net_29            = 4'h0;
assign OE_DATA_124_const_net_29            = 4'h0;
assign OE_DATA_125_const_net_29            = 4'h0;
assign OE_DATA_126_const_net_29            = 4'h0;
assign OE_DATA_127_const_net_29            = 4'h0;
assign CDR_CLK_B_SEL_const_net_3           = 11'h000;
assign FIFO_WR_PTR_const_net_21            = 3'h0;
assign FIFO_RD_PTR_const_net_21            = 3'h0;
assign EYE_MONITOR_LANE_WIDTH_const_net_24 = 3'h0;
assign TX_DATA_1_const_net_24              = 8'h00;
assign TX_DATA_2_const_net_26              = 8'h00;
assign TX_DATA_3_const_net_26              = 8'h00;
assign TX_DATA_4_const_net_26              = 8'h00;
assign TX_DATA_5_const_net_26              = 8'h00;
assign TX_DATA_6_const_net_26              = 8'h00;
assign TX_DATA_7_const_net_26              = 8'h00;
assign TX_DATA_8_const_net_29              = 8'h00;
assign TX_DATA_9_const_net_29              = 8'h00;
assign TX_DATA_10_const_net_29             = 8'h00;
assign TX_DATA_11_const_net_29             = 8'h00;
assign TX_DATA_12_const_net_30             = 8'h00;
assign TX_DATA_13_const_net_30             = 8'h00;
assign TX_DATA_14_const_net_30             = 8'h00;
assign TX_DATA_15_const_net_30             = 8'h00;
assign TX_DATA_16_const_net_30             = 8'h00;
assign TX_DATA_17_const_net_30             = 8'h00;
assign TX_DATA_18_const_net_30             = 8'h00;
assign TX_DATA_19_const_net_30             = 8'h00;
assign TX_DATA_20_const_net_30             = 8'h00;
assign TX_DATA_21_const_net_30             = 8'h00;
assign TX_DATA_22_const_net_30             = 8'h00;
assign TX_DATA_23_const_net_30             = 8'h00;
assign TX_DATA_24_const_net_30             = 8'h00;
assign TX_DATA_25_const_net_30             = 8'h00;
assign TX_DATA_26_const_net_30             = 8'h00;
assign TX_DATA_27_const_net_30             = 8'h00;
assign TX_DATA_28_const_net_30             = 8'h00;
assign TX_DATA_29_const_net_30             = 8'h00;
assign TX_DATA_30_const_net_30             = 8'h00;
assign TX_DATA_31_const_net_30             = 8'h00;
assign TX_DATA_32_const_net_30             = 8'h00;
assign TX_DATA_33_const_net_30             = 8'h00;
assign TX_DATA_34_const_net_30             = 8'h00;
assign TX_DATA_35_const_net_30             = 8'h00;
assign TX_DATA_36_const_net_30             = 8'h00;
assign TX_DATA_37_const_net_30             = 8'h00;
assign TX_DATA_38_const_net_30             = 8'h00;
assign TX_DATA_39_const_net_30             = 8'h00;
assign TX_DATA_40_const_net_30             = 8'h00;
assign TX_DATA_41_const_net_30             = 8'h00;
assign TX_DATA_42_const_net_30             = 8'h00;
assign TX_DATA_43_const_net_30             = 8'h00;
assign TX_DATA_44_const_net_30             = 8'h00;
assign TX_DATA_45_const_net_30             = 8'h00;
assign TX_DATA_46_const_net_30             = 8'h00;
assign TX_DATA_47_const_net_30             = 8'h00;
assign TX_DATA_48_const_net_30             = 8'h00;
assign TX_DATA_49_const_net_30             = 8'h00;
assign TX_DATA_50_const_net_30             = 8'h00;
assign TX_DATA_51_const_net_30             = 8'h00;
assign TX_DATA_52_const_net_30             = 8'h00;
assign TX_DATA_53_const_net_30             = 8'h00;
assign TX_DATA_54_const_net_30             = 8'h00;
assign TX_DATA_55_const_net_30             = 8'h00;
assign TX_DATA_56_const_net_30             = 8'h00;
assign TX_DATA_57_const_net_30             = 8'h00;
assign TX_DATA_58_const_net_30             = 8'h00;
assign TX_DATA_59_const_net_30             = 8'h00;
assign TX_DATA_60_const_net_30             = 8'h00;
assign TX_DATA_61_const_net_30             = 8'h00;
assign TX_DATA_62_const_net_30             = 8'h00;
assign TX_DATA_63_const_net_30             = 8'h00;
assign TX_DATA_64_const_net_30             = 8'h00;
assign TX_DATA_65_const_net_30             = 8'h00;
assign TX_DATA_66_const_net_30             = 8'h00;
assign TX_DATA_67_const_net_30             = 8'h00;
assign TX_DATA_68_const_net_30             = 8'h00;
assign TX_DATA_69_const_net_30             = 8'h00;
assign TX_DATA_70_const_net_30             = 8'h00;
assign TX_DATA_71_const_net_30             = 8'h00;
assign TX_DATA_72_const_net_30             = 8'h00;
assign TX_DATA_73_const_net_30             = 8'h00;
assign TX_DATA_74_const_net_30             = 8'h00;
assign TX_DATA_75_const_net_30             = 8'h00;
assign TX_DATA_76_const_net_30             = 8'h00;
assign TX_DATA_77_const_net_30             = 8'h00;
assign TX_DATA_78_const_net_30             = 8'h00;
assign TX_DATA_79_const_net_30             = 8'h00;
assign TX_DATA_80_const_net_30             = 8'h00;
assign TX_DATA_81_const_net_30             = 8'h00;
assign TX_DATA_82_const_net_30             = 8'h00;
assign TX_DATA_83_const_net_30             = 8'h00;
assign TX_DATA_84_const_net_30             = 8'h00;
assign TX_DATA_85_const_net_30             = 8'h00;
assign TX_DATA_86_const_net_30             = 8'h00;
assign TX_DATA_87_const_net_30             = 8'h00;
assign TX_DATA_88_const_net_30             = 8'h00;
assign TX_DATA_89_const_net_30             = 8'h00;
assign TX_DATA_90_const_net_30             = 8'h00;
assign TX_DATA_91_const_net_30             = 8'h00;
assign TX_DATA_92_const_net_30             = 8'h00;
assign TX_DATA_93_const_net_30             = 8'h00;
assign TX_DATA_94_const_net_30             = 8'h00;
assign TX_DATA_95_const_net_30             = 8'h00;
assign TX_DATA_96_const_net_30             = 8'h00;
assign TX_DATA_97_const_net_30             = 8'h00;
assign TX_DATA_98_const_net_30             = 8'h00;
assign TX_DATA_99_const_net_30             = 8'h00;
assign TX_DATA_100_const_net_30            = 8'h00;
assign TX_DATA_101_const_net_30            = 8'h00;
assign TX_DATA_102_const_net_30            = 8'h00;
assign TX_DATA_103_const_net_30            = 8'h00;
assign TX_DATA_104_const_net_30            = 8'h00;
assign TX_DATA_105_const_net_30            = 8'h00;
assign TX_DATA_106_const_net_30            = 8'h00;
assign TX_DATA_107_const_net_30            = 8'h00;
assign TX_DATA_108_const_net_30            = 8'h00;
assign TX_DATA_109_const_net_30            = 8'h00;
assign TX_DATA_110_const_net_30            = 8'h00;
assign TX_DATA_111_const_net_30            = 8'h00;
assign TX_DATA_112_const_net_30            = 8'h00;
assign TX_DATA_113_const_net_30            = 8'h00;
assign TX_DATA_114_const_net_30            = 8'h00;
assign TX_DATA_115_const_net_30            = 8'h00;
assign TX_DATA_116_const_net_30            = 8'h00;
assign TX_DATA_117_const_net_30            = 8'h00;
assign TX_DATA_118_const_net_30            = 8'h00;
assign TX_DATA_119_const_net_30            = 8'h00;
assign TX_DATA_120_const_net_30            = 8'h00;
assign TX_DATA_121_const_net_30            = 8'h00;
assign TX_DATA_122_const_net_30            = 8'h00;
assign TX_DATA_123_const_net_30            = 8'h00;
assign TX_DATA_124_const_net_30            = 8'h00;
assign TX_DATA_125_const_net_30            = 8'h00;
assign TX_DATA_126_const_net_30            = 8'h00;
assign TX_DATA_127_const_net_30            = 8'h00;
assign OE_DATA_1_const_net_27              = 4'h0;
assign OE_DATA_2_const_net_27              = 4'h0;
assign OE_DATA_3_const_net_27              = 4'h0;
assign OE_DATA_4_const_net_27              = 4'h0;
assign OE_DATA_5_const_net_27              = 4'h0;
assign OE_DATA_6_const_net_27              = 4'h0;
assign OE_DATA_7_const_net_27              = 4'h0;
assign OE_DATA_8_const_net_30              = 4'h0;
assign OE_DATA_9_const_net_30              = 4'h0;
assign OE_DATA_10_const_net_30             = 4'h0;
assign OE_DATA_11_const_net_30             = 4'h0;
assign OE_DATA_12_const_net_30             = 4'h0;
assign OE_DATA_13_const_net_30             = 4'h0;
assign OE_DATA_14_const_net_30             = 4'h0;
assign OE_DATA_15_const_net_30             = 4'h0;
assign OE_DATA_16_const_net_30             = 4'h0;
assign OE_DATA_17_const_net_30             = 4'h0;
assign OE_DATA_18_const_net_30             = 4'h0;
assign OE_DATA_19_const_net_30             = 4'h0;
assign OE_DATA_20_const_net_30             = 4'h0;
assign OE_DATA_21_const_net_30             = 4'h0;
assign OE_DATA_22_const_net_30             = 4'h0;
assign OE_DATA_23_const_net_30             = 4'h0;
assign OE_DATA_24_const_net_30             = 4'h0;
assign OE_DATA_25_const_net_30             = 4'h0;
assign OE_DATA_26_const_net_30             = 4'h0;
assign OE_DATA_27_const_net_30             = 4'h0;
assign OE_DATA_28_const_net_30             = 4'h0;
assign OE_DATA_29_const_net_30             = 4'h0;
assign OE_DATA_30_const_net_30             = 4'h0;
assign OE_DATA_31_const_net_30             = 4'h0;
assign OE_DATA_32_const_net_30             = 4'h0;
assign OE_DATA_33_const_net_30             = 4'h0;
assign OE_DATA_34_const_net_30             = 4'h0;
assign OE_DATA_35_const_net_30             = 4'h0;
assign OE_DATA_36_const_net_30             = 4'h0;
assign OE_DATA_37_const_net_30             = 4'h0;
assign OE_DATA_38_const_net_30             = 4'h0;
assign OE_DATA_39_const_net_30             = 4'h0;
assign OE_DATA_40_const_net_30             = 4'h0;
assign OE_DATA_41_const_net_30             = 4'h0;
assign OE_DATA_42_const_net_30             = 4'h0;
assign OE_DATA_43_const_net_30             = 4'h0;
assign OE_DATA_44_const_net_30             = 4'h0;
assign OE_DATA_45_const_net_30             = 4'h0;
assign OE_DATA_46_const_net_30             = 4'h0;
assign OE_DATA_47_const_net_30             = 4'h0;
assign OE_DATA_48_const_net_30             = 4'h0;
assign OE_DATA_49_const_net_30             = 4'h0;
assign OE_DATA_50_const_net_30             = 4'h0;
assign OE_DATA_51_const_net_30             = 4'h0;
assign OE_DATA_52_const_net_30             = 4'h0;
assign OE_DATA_53_const_net_30             = 4'h0;
assign OE_DATA_54_const_net_30             = 4'h0;
assign OE_DATA_55_const_net_30             = 4'h0;
assign OE_DATA_56_const_net_30             = 4'h0;
assign OE_DATA_57_const_net_30             = 4'h0;
assign OE_DATA_58_const_net_30             = 4'h0;
assign OE_DATA_59_const_net_30             = 4'h0;
assign OE_DATA_60_const_net_30             = 4'h0;
assign OE_DATA_61_const_net_30             = 4'h0;
assign OE_DATA_62_const_net_30             = 4'h0;
assign OE_DATA_63_const_net_30             = 4'h0;
assign OE_DATA_64_const_net_30             = 4'h0;
assign OE_DATA_65_const_net_30             = 4'h0;
assign OE_DATA_66_const_net_30             = 4'h0;
assign OE_DATA_67_const_net_30             = 4'h0;
assign OE_DATA_68_const_net_30             = 4'h0;
assign OE_DATA_69_const_net_30             = 4'h0;
assign OE_DATA_70_const_net_30             = 4'h0;
assign OE_DATA_71_const_net_30             = 4'h0;
assign OE_DATA_72_const_net_30             = 4'h0;
assign OE_DATA_73_const_net_30             = 4'h0;
assign OE_DATA_74_const_net_30             = 4'h0;
assign OE_DATA_75_const_net_30             = 4'h0;
assign OE_DATA_76_const_net_30             = 4'h0;
assign OE_DATA_77_const_net_30             = 4'h0;
assign OE_DATA_78_const_net_30             = 4'h0;
assign OE_DATA_79_const_net_30             = 4'h0;
assign OE_DATA_80_const_net_30             = 4'h0;
assign OE_DATA_81_const_net_30             = 4'h0;
assign OE_DATA_82_const_net_30             = 4'h0;
assign OE_DATA_83_const_net_30             = 4'h0;
assign OE_DATA_84_const_net_30             = 4'h0;
assign OE_DATA_85_const_net_30             = 4'h0;
assign OE_DATA_86_const_net_30             = 4'h0;
assign OE_DATA_87_const_net_30             = 4'h0;
assign OE_DATA_88_const_net_30             = 4'h0;
assign OE_DATA_89_const_net_30             = 4'h0;
assign OE_DATA_90_const_net_30             = 4'h0;
assign OE_DATA_91_const_net_30             = 4'h0;
assign OE_DATA_92_const_net_30             = 4'h0;
assign OE_DATA_93_const_net_30             = 4'h0;
assign OE_DATA_94_const_net_30             = 4'h0;
assign OE_DATA_95_const_net_30             = 4'h0;
assign OE_DATA_96_const_net_30             = 4'h0;
assign OE_DATA_97_const_net_30             = 4'h0;
assign OE_DATA_98_const_net_30             = 4'h0;
assign OE_DATA_99_const_net_30             = 4'h0;
assign OE_DATA_100_const_net_30            = 4'h0;
assign OE_DATA_101_const_net_30            = 4'h0;
assign OE_DATA_102_const_net_30            = 4'h0;
assign OE_DATA_103_const_net_30            = 4'h0;
assign OE_DATA_104_const_net_30            = 4'h0;
assign OE_DATA_105_const_net_30            = 4'h0;
assign OE_DATA_106_const_net_30            = 4'h0;
assign OE_DATA_107_const_net_30            = 4'h0;
assign OE_DATA_108_const_net_30            = 4'h0;
assign OE_DATA_109_const_net_30            = 4'h0;
assign OE_DATA_110_const_net_30            = 4'h0;
assign OE_DATA_111_const_net_30            = 4'h0;
assign OE_DATA_112_const_net_30            = 4'h0;
assign OE_DATA_113_const_net_30            = 4'h0;
assign OE_DATA_114_const_net_30            = 4'h0;
assign OE_DATA_115_const_net_30            = 4'h0;
assign OE_DATA_116_const_net_30            = 4'h0;
assign OE_DATA_117_const_net_30            = 4'h0;
assign OE_DATA_118_const_net_30            = 4'h0;
assign OE_DATA_119_const_net_30            = 4'h0;
assign OE_DATA_120_const_net_30            = 4'h0;
assign OE_DATA_121_const_net_30            = 4'h0;
assign OE_DATA_122_const_net_30            = 4'h0;
assign OE_DATA_123_const_net_30            = 4'h0;
assign OE_DATA_124_const_net_30            = 4'h0;
assign OE_DATA_125_const_net_30            = 4'h0;
assign OE_DATA_126_const_net_30            = 4'h0;
assign OE_DATA_127_const_net_30            = 4'h0;
assign TX_DATA_8_const_net_30              = 8'h00;
assign TX_DATA_9_const_net_30              = 8'h00;
assign TX_DATA_10_const_net_30             = 8'h00;
assign TX_DATA_11_const_net_30             = 8'h00;
assign TX_DATA_12_const_net_31             = 8'h00;
assign TX_DATA_13_const_net_31             = 8'h00;
assign TX_DATA_14_const_net_31             = 8'h00;
assign TX_DATA_15_const_net_31             = 8'h00;
assign TX_DATA_16_const_net_31             = 8'h00;
assign TX_DATA_17_const_net_31             = 8'h00;
assign TX_DATA_18_const_net_31             = 8'h00;
assign TX_DATA_19_const_net_31             = 8'h00;
assign TX_DATA_20_const_net_31             = 8'h00;
assign TX_DATA_21_const_net_31             = 8'h00;
assign TX_DATA_22_const_net_31             = 8'h00;
assign TX_DATA_23_const_net_31             = 8'h00;
assign TX_DATA_24_const_net_31             = 8'h00;
assign TX_DATA_25_const_net_31             = 8'h00;
assign TX_DATA_26_const_net_31             = 8'h00;
assign TX_DATA_27_const_net_31             = 8'h00;
assign TX_DATA_28_const_net_31             = 8'h00;
assign TX_DATA_29_const_net_31             = 8'h00;
assign TX_DATA_30_const_net_31             = 8'h00;
assign TX_DATA_31_const_net_31             = 8'h00;
assign TX_DATA_32_const_net_31             = 8'h00;
assign TX_DATA_33_const_net_31             = 8'h00;
assign TX_DATA_34_const_net_31             = 8'h00;
assign TX_DATA_35_const_net_31             = 8'h00;
assign TX_DATA_36_const_net_31             = 8'h00;
assign TX_DATA_37_const_net_31             = 8'h00;
assign TX_DATA_38_const_net_31             = 8'h00;
assign TX_DATA_39_const_net_31             = 8'h00;
assign TX_DATA_40_const_net_31             = 8'h00;
assign TX_DATA_41_const_net_31             = 8'h00;
assign TX_DATA_42_const_net_31             = 8'h00;
assign TX_DATA_43_const_net_31             = 8'h00;
assign TX_DATA_44_const_net_31             = 8'h00;
assign TX_DATA_45_const_net_31             = 8'h00;
assign TX_DATA_46_const_net_31             = 8'h00;
assign TX_DATA_47_const_net_31             = 8'h00;
assign TX_DATA_48_const_net_31             = 8'h00;
assign TX_DATA_49_const_net_31             = 8'h00;
assign TX_DATA_50_const_net_31             = 8'h00;
assign TX_DATA_51_const_net_31             = 8'h00;
assign TX_DATA_52_const_net_31             = 8'h00;
assign TX_DATA_53_const_net_31             = 8'h00;
assign TX_DATA_54_const_net_31             = 8'h00;
assign TX_DATA_55_const_net_31             = 8'h00;
assign TX_DATA_56_const_net_31             = 8'h00;
assign TX_DATA_57_const_net_31             = 8'h00;
assign TX_DATA_58_const_net_31             = 8'h00;
assign TX_DATA_59_const_net_31             = 8'h00;
assign TX_DATA_60_const_net_31             = 8'h00;
assign TX_DATA_61_const_net_31             = 8'h00;
assign TX_DATA_62_const_net_31             = 8'h00;
assign TX_DATA_63_const_net_31             = 8'h00;
assign TX_DATA_64_const_net_31             = 8'h00;
assign TX_DATA_65_const_net_31             = 8'h00;
assign TX_DATA_66_const_net_31             = 8'h00;
assign TX_DATA_67_const_net_31             = 8'h00;
assign TX_DATA_68_const_net_31             = 8'h00;
assign TX_DATA_69_const_net_31             = 8'h00;
assign TX_DATA_70_const_net_31             = 8'h00;
assign TX_DATA_71_const_net_31             = 8'h00;
assign TX_DATA_72_const_net_31             = 8'h00;
assign TX_DATA_73_const_net_31             = 8'h00;
assign TX_DATA_74_const_net_31             = 8'h00;
assign TX_DATA_75_const_net_31             = 8'h00;
assign TX_DATA_76_const_net_31             = 8'h00;
assign TX_DATA_77_const_net_31             = 8'h00;
assign TX_DATA_78_const_net_31             = 8'h00;
assign TX_DATA_79_const_net_31             = 8'h00;
assign TX_DATA_80_const_net_31             = 8'h00;
assign TX_DATA_81_const_net_31             = 8'h00;
assign TX_DATA_82_const_net_31             = 8'h00;
assign TX_DATA_83_const_net_31             = 8'h00;
assign TX_DATA_84_const_net_31             = 8'h00;
assign TX_DATA_85_const_net_31             = 8'h00;
assign TX_DATA_86_const_net_31             = 8'h00;
assign TX_DATA_87_const_net_31             = 8'h00;
assign TX_DATA_88_const_net_31             = 8'h00;
assign TX_DATA_89_const_net_31             = 8'h00;
assign TX_DATA_90_const_net_31             = 8'h00;
assign TX_DATA_91_const_net_31             = 8'h00;
assign TX_DATA_92_const_net_31             = 8'h00;
assign TX_DATA_93_const_net_31             = 8'h00;
assign TX_DATA_94_const_net_31             = 8'h00;
assign TX_DATA_95_const_net_31             = 8'h00;
assign TX_DATA_96_const_net_31             = 8'h00;
assign TX_DATA_97_const_net_31             = 8'h00;
assign TX_DATA_98_const_net_31             = 8'h00;
assign TX_DATA_99_const_net_31             = 8'h00;
assign TX_DATA_100_const_net_31            = 8'h00;
assign TX_DATA_101_const_net_31            = 8'h00;
assign TX_DATA_102_const_net_31            = 8'h00;
assign TX_DATA_103_const_net_31            = 8'h00;
assign TX_DATA_104_const_net_31            = 8'h00;
assign TX_DATA_105_const_net_31            = 8'h00;
assign TX_DATA_106_const_net_31            = 8'h00;
assign TX_DATA_107_const_net_31            = 8'h00;
assign TX_DATA_108_const_net_31            = 8'h00;
assign TX_DATA_109_const_net_31            = 8'h00;
assign TX_DATA_110_const_net_31            = 8'h00;
assign TX_DATA_111_const_net_31            = 8'h00;
assign TX_DATA_112_const_net_31            = 8'h00;
assign TX_DATA_113_const_net_31            = 8'h00;
assign TX_DATA_114_const_net_31            = 8'h00;
assign TX_DATA_115_const_net_31            = 8'h00;
assign TX_DATA_116_const_net_31            = 8'h00;
assign TX_DATA_117_const_net_31            = 8'h00;
assign TX_DATA_118_const_net_31            = 8'h00;
assign TX_DATA_119_const_net_31            = 8'h00;
assign TX_DATA_120_const_net_31            = 8'h00;
assign TX_DATA_121_const_net_31            = 8'h00;
assign TX_DATA_122_const_net_31            = 8'h00;
assign TX_DATA_123_const_net_31            = 8'h00;
assign TX_DATA_124_const_net_31            = 8'h00;
assign TX_DATA_125_const_net_31            = 8'h00;
assign TX_DATA_126_const_net_31            = 8'h00;
assign TX_DATA_127_const_net_31            = 8'h00;
assign OE_DATA_8_const_net_31              = 4'h0;
assign OE_DATA_9_const_net_31              = 4'h0;
assign OE_DATA_10_const_net_31             = 4'h0;
assign OE_DATA_11_const_net_31             = 4'h0;
assign OE_DATA_12_const_net_31             = 4'h0;
assign OE_DATA_13_const_net_31             = 4'h0;
assign OE_DATA_14_const_net_31             = 4'h0;
assign OE_DATA_15_const_net_31             = 4'h0;
assign OE_DATA_16_const_net_31             = 4'h0;
assign OE_DATA_17_const_net_31             = 4'h0;
assign OE_DATA_18_const_net_31             = 4'h0;
assign OE_DATA_19_const_net_31             = 4'h0;
assign OE_DATA_20_const_net_31             = 4'h0;
assign OE_DATA_21_const_net_31             = 4'h0;
assign OE_DATA_22_const_net_31             = 4'h0;
assign OE_DATA_23_const_net_31             = 4'h0;
assign OE_DATA_24_const_net_31             = 4'h0;
assign OE_DATA_25_const_net_31             = 4'h0;
assign OE_DATA_26_const_net_31             = 4'h0;
assign OE_DATA_27_const_net_31             = 4'h0;
assign OE_DATA_28_const_net_31             = 4'h0;
assign OE_DATA_29_const_net_31             = 4'h0;
assign OE_DATA_30_const_net_31             = 4'h0;
assign OE_DATA_31_const_net_31             = 4'h0;
assign OE_DATA_32_const_net_31             = 4'h0;
assign OE_DATA_33_const_net_31             = 4'h0;
assign OE_DATA_34_const_net_31             = 4'h0;
assign OE_DATA_35_const_net_31             = 4'h0;
assign OE_DATA_36_const_net_31             = 4'h0;
assign OE_DATA_37_const_net_31             = 4'h0;
assign OE_DATA_38_const_net_31             = 4'h0;
assign OE_DATA_39_const_net_31             = 4'h0;
assign OE_DATA_40_const_net_31             = 4'h0;
assign OE_DATA_41_const_net_31             = 4'h0;
assign OE_DATA_42_const_net_31             = 4'h0;
assign OE_DATA_43_const_net_31             = 4'h0;
assign OE_DATA_44_const_net_31             = 4'h0;
assign OE_DATA_45_const_net_31             = 4'h0;
assign OE_DATA_46_const_net_31             = 4'h0;
assign OE_DATA_47_const_net_31             = 4'h0;
assign OE_DATA_48_const_net_31             = 4'h0;
assign OE_DATA_49_const_net_31             = 4'h0;
assign OE_DATA_50_const_net_31             = 4'h0;
assign OE_DATA_51_const_net_31             = 4'h0;
assign OE_DATA_52_const_net_31             = 4'h0;
assign OE_DATA_53_const_net_31             = 4'h0;
assign OE_DATA_54_const_net_31             = 4'h0;
assign OE_DATA_55_const_net_31             = 4'h0;
assign OE_DATA_56_const_net_31             = 4'h0;
assign OE_DATA_57_const_net_31             = 4'h0;
assign OE_DATA_58_const_net_31             = 4'h0;
assign OE_DATA_59_const_net_31             = 4'h0;
assign OE_DATA_60_const_net_31             = 4'h0;
assign OE_DATA_61_const_net_31             = 4'h0;
assign OE_DATA_62_const_net_31             = 4'h0;
assign OE_DATA_63_const_net_31             = 4'h0;
assign OE_DATA_64_const_net_31             = 4'h0;
assign OE_DATA_65_const_net_31             = 4'h0;
assign OE_DATA_66_const_net_31             = 4'h0;
assign OE_DATA_67_const_net_31             = 4'h0;
assign OE_DATA_68_const_net_31             = 4'h0;
assign OE_DATA_69_const_net_31             = 4'h0;
assign OE_DATA_70_const_net_31             = 4'h0;
assign OE_DATA_71_const_net_31             = 4'h0;
assign OE_DATA_72_const_net_31             = 4'h0;
assign OE_DATA_73_const_net_31             = 4'h0;
assign OE_DATA_74_const_net_31             = 4'h0;
assign OE_DATA_75_const_net_31             = 4'h0;
assign OE_DATA_76_const_net_31             = 4'h0;
assign OE_DATA_77_const_net_31             = 4'h0;
assign OE_DATA_78_const_net_31             = 4'h0;
assign OE_DATA_79_const_net_31             = 4'h0;
assign OE_DATA_80_const_net_31             = 4'h0;
assign OE_DATA_81_const_net_31             = 4'h0;
assign OE_DATA_82_const_net_31             = 4'h0;
assign OE_DATA_83_const_net_31             = 4'h0;
assign OE_DATA_84_const_net_31             = 4'h0;
assign OE_DATA_85_const_net_31             = 4'h0;
assign OE_DATA_86_const_net_31             = 4'h0;
assign OE_DATA_87_const_net_31             = 4'h0;
assign OE_DATA_88_const_net_31             = 4'h0;
assign OE_DATA_89_const_net_31             = 4'h0;
assign OE_DATA_90_const_net_31             = 4'h0;
assign OE_DATA_91_const_net_31             = 4'h0;
assign OE_DATA_92_const_net_31             = 4'h0;
assign OE_DATA_93_const_net_31             = 4'h0;
assign OE_DATA_94_const_net_31             = 4'h0;
assign OE_DATA_95_const_net_31             = 4'h0;
assign OE_DATA_96_const_net_31             = 4'h0;
assign OE_DATA_97_const_net_31             = 4'h0;
assign OE_DATA_98_const_net_31             = 4'h0;
assign OE_DATA_99_const_net_31             = 4'h0;
assign OE_DATA_100_const_net_31            = 4'h0;
assign OE_DATA_101_const_net_31            = 4'h0;
assign OE_DATA_102_const_net_31            = 4'h0;
assign OE_DATA_103_const_net_31            = 4'h0;
assign OE_DATA_104_const_net_31            = 4'h0;
assign OE_DATA_105_const_net_31            = 4'h0;
assign OE_DATA_106_const_net_31            = 4'h0;
assign OE_DATA_107_const_net_31            = 4'h0;
assign OE_DATA_108_const_net_31            = 4'h0;
assign OE_DATA_109_const_net_31            = 4'h0;
assign OE_DATA_110_const_net_31            = 4'h0;
assign OE_DATA_111_const_net_31            = 4'h0;
assign OE_DATA_112_const_net_31            = 4'h0;
assign OE_DATA_113_const_net_31            = 4'h0;
assign OE_DATA_114_const_net_31            = 4'h0;
assign OE_DATA_115_const_net_31            = 4'h0;
assign OE_DATA_116_const_net_31            = 4'h0;
assign OE_DATA_117_const_net_31            = 4'h0;
assign OE_DATA_118_const_net_31            = 4'h0;
assign OE_DATA_119_const_net_31            = 4'h0;
assign OE_DATA_120_const_net_31            = 4'h0;
assign OE_DATA_121_const_net_31            = 4'h0;
assign OE_DATA_122_const_net_31            = 4'h0;
assign OE_DATA_123_const_net_31            = 4'h0;
assign OE_DATA_124_const_net_31            = 4'h0;
assign OE_DATA_125_const_net_31            = 4'h0;
assign OE_DATA_126_const_net_31            = 4'h0;
assign OE_DATA_127_const_net_31            = 4'h0;
assign PAD_I_const_net_6                   = 8'h00;
assign PAD_N_const_net_6                   = 8'h00;
assign PAD_I_N_const_net_6                 = 8'h00;
assign TX_DATA_1_const_net_25              = 8'h00;
assign TX_DATA_2_const_net_27              = 8'h00;
assign TX_DATA_3_const_net_27              = 8'h00;
assign TX_DATA_4_const_net_27              = 8'h00;
assign TX_DATA_5_const_net_27              = 8'h00;
assign TX_DATA_6_const_net_27              = 8'h00;
assign TX_DATA_7_const_net_27              = 8'h00;
assign TX_DATA_8_const_net_31              = 8'h00;
assign TX_DATA_9_const_net_31              = 8'h00;
assign TX_DATA_10_const_net_31             = 8'h00;
assign TX_DATA_11_const_net_31             = 8'h00;
assign TX_DATA_12_const_net_32             = 8'h00;
assign TX_DATA_13_const_net_32             = 8'h00;
assign TX_DATA_14_const_net_32             = 8'h00;
assign TX_DATA_15_const_net_32             = 8'h00;
assign TX_DATA_16_const_net_32             = 8'h00;
assign TX_DATA_17_const_net_32             = 8'h00;
assign TX_DATA_18_const_net_32             = 8'h00;
assign TX_DATA_19_const_net_32             = 8'h00;
assign TX_DATA_20_const_net_32             = 8'h00;
assign TX_DATA_21_const_net_32             = 8'h00;
assign TX_DATA_22_const_net_32             = 8'h00;
assign TX_DATA_23_const_net_32             = 8'h00;
assign TX_DATA_24_const_net_32             = 8'h00;
assign TX_DATA_25_const_net_32             = 8'h00;
assign TX_DATA_26_const_net_32             = 8'h00;
assign TX_DATA_27_const_net_32             = 8'h00;
assign TX_DATA_28_const_net_32             = 8'h00;
assign TX_DATA_29_const_net_32             = 8'h00;
assign TX_DATA_30_const_net_32             = 8'h00;
assign TX_DATA_31_const_net_32             = 8'h00;
assign TX_DATA_32_const_net_32             = 8'h00;
assign TX_DATA_33_const_net_32             = 8'h00;
assign TX_DATA_34_const_net_32             = 8'h00;
assign TX_DATA_35_const_net_32             = 8'h00;
assign TX_DATA_36_const_net_32             = 8'h00;
assign TX_DATA_37_const_net_32             = 8'h00;
assign TX_DATA_38_const_net_32             = 8'h00;
assign TX_DATA_39_const_net_32             = 8'h00;
assign TX_DATA_40_const_net_32             = 8'h00;
assign TX_DATA_41_const_net_32             = 8'h00;
assign TX_DATA_42_const_net_32             = 8'h00;
assign TX_DATA_43_const_net_32             = 8'h00;
assign TX_DATA_44_const_net_32             = 8'h00;
assign TX_DATA_45_const_net_32             = 8'h00;
assign TX_DATA_46_const_net_32             = 8'h00;
assign TX_DATA_47_const_net_32             = 8'h00;
assign TX_DATA_48_const_net_32             = 8'h00;
assign TX_DATA_49_const_net_32             = 8'h00;
assign TX_DATA_50_const_net_32             = 8'h00;
assign TX_DATA_51_const_net_32             = 8'h00;
assign TX_DATA_52_const_net_32             = 8'h00;
assign TX_DATA_53_const_net_32             = 8'h00;
assign TX_DATA_54_const_net_32             = 8'h00;
assign TX_DATA_55_const_net_32             = 8'h00;
assign TX_DATA_56_const_net_32             = 8'h00;
assign TX_DATA_57_const_net_32             = 8'h00;
assign TX_DATA_58_const_net_32             = 8'h00;
assign TX_DATA_59_const_net_32             = 8'h00;
assign TX_DATA_60_const_net_32             = 8'h00;
assign TX_DATA_61_const_net_32             = 8'h00;
assign TX_DATA_62_const_net_32             = 8'h00;
assign TX_DATA_63_const_net_32             = 8'h00;
assign TX_DATA_64_const_net_32             = 8'h00;
assign TX_DATA_65_const_net_32             = 8'h00;
assign TX_DATA_66_const_net_32             = 8'h00;
assign TX_DATA_67_const_net_32             = 8'h00;
assign TX_DATA_68_const_net_32             = 8'h00;
assign TX_DATA_69_const_net_32             = 8'h00;
assign TX_DATA_70_const_net_32             = 8'h00;
assign TX_DATA_71_const_net_32             = 8'h00;
assign TX_DATA_72_const_net_32             = 8'h00;
assign TX_DATA_73_const_net_32             = 8'h00;
assign TX_DATA_74_const_net_32             = 8'h00;
assign TX_DATA_75_const_net_32             = 8'h00;
assign TX_DATA_76_const_net_32             = 8'h00;
assign TX_DATA_77_const_net_32             = 8'h00;
assign TX_DATA_78_const_net_32             = 8'h00;
assign TX_DATA_79_const_net_32             = 8'h00;
assign TX_DATA_80_const_net_32             = 8'h00;
assign TX_DATA_81_const_net_32             = 8'h00;
assign TX_DATA_82_const_net_32             = 8'h00;
assign TX_DATA_83_const_net_32             = 8'h00;
assign TX_DATA_84_const_net_32             = 8'h00;
assign TX_DATA_85_const_net_32             = 8'h00;
assign TX_DATA_86_const_net_32             = 8'h00;
assign TX_DATA_87_const_net_32             = 8'h00;
assign TX_DATA_88_const_net_32             = 8'h00;
assign TX_DATA_89_const_net_32             = 8'h00;
assign TX_DATA_90_const_net_32             = 8'h00;
assign TX_DATA_91_const_net_32             = 8'h00;
assign TX_DATA_92_const_net_32             = 8'h00;
assign TX_DATA_93_const_net_32             = 8'h00;
assign TX_DATA_94_const_net_32             = 8'h00;
assign TX_DATA_95_const_net_32             = 8'h00;
assign TX_DATA_96_const_net_32             = 8'h00;
assign TX_DATA_97_const_net_32             = 8'h00;
assign TX_DATA_98_const_net_32             = 8'h00;
assign TX_DATA_99_const_net_32             = 8'h00;
assign TX_DATA_100_const_net_32            = 8'h00;
assign TX_DATA_101_const_net_32            = 8'h00;
assign TX_DATA_102_const_net_32            = 8'h00;
assign TX_DATA_103_const_net_32            = 8'h00;
assign TX_DATA_104_const_net_32            = 8'h00;
assign TX_DATA_105_const_net_32            = 8'h00;
assign TX_DATA_106_const_net_32            = 8'h00;
assign TX_DATA_107_const_net_32            = 8'h00;
assign TX_DATA_108_const_net_32            = 8'h00;
assign TX_DATA_109_const_net_32            = 8'h00;
assign TX_DATA_110_const_net_32            = 8'h00;
assign TX_DATA_111_const_net_32            = 8'h00;
assign TX_DATA_112_const_net_32            = 8'h00;
assign TX_DATA_113_const_net_32            = 8'h00;
assign TX_DATA_114_const_net_32            = 8'h00;
assign TX_DATA_115_const_net_32            = 8'h00;
assign TX_DATA_116_const_net_32            = 8'h00;
assign TX_DATA_117_const_net_32            = 8'h00;
assign TX_DATA_118_const_net_32            = 8'h00;
assign TX_DATA_119_const_net_32            = 8'h00;
assign TX_DATA_120_const_net_32            = 8'h00;
assign TX_DATA_121_const_net_32            = 8'h00;
assign TX_DATA_122_const_net_32            = 8'h00;
assign TX_DATA_123_const_net_32            = 8'h00;
assign TX_DATA_124_const_net_32            = 8'h00;
assign TX_DATA_125_const_net_32            = 8'h00;
assign TX_DATA_126_const_net_32            = 8'h00;
assign TX_DATA_127_const_net_32            = 8'h00;
assign OE_DATA_1_const_net_28              = 4'h0;
assign OE_DATA_2_const_net_28              = 4'h0;
assign OE_DATA_3_const_net_28              = 4'h0;
assign OE_DATA_4_const_net_28              = 4'h0;
assign OE_DATA_5_const_net_28              = 4'h0;
assign OE_DATA_6_const_net_28              = 4'h0;
assign OE_DATA_7_const_net_28              = 4'h0;
assign OE_DATA_8_const_net_32              = 4'h0;
assign OE_DATA_9_const_net_32              = 4'h0;
assign OE_DATA_10_const_net_32             = 4'h0;
assign OE_DATA_11_const_net_32             = 4'h0;
assign OE_DATA_12_const_net_32             = 4'h0;
assign OE_DATA_13_const_net_32             = 4'h0;
assign OE_DATA_14_const_net_32             = 4'h0;
assign OE_DATA_15_const_net_32             = 4'h0;
assign OE_DATA_16_const_net_32             = 4'h0;
assign OE_DATA_17_const_net_32             = 4'h0;
assign OE_DATA_18_const_net_32             = 4'h0;
assign OE_DATA_19_const_net_32             = 4'h0;
assign OE_DATA_20_const_net_32             = 4'h0;
assign OE_DATA_21_const_net_32             = 4'h0;
assign OE_DATA_22_const_net_32             = 4'h0;
assign OE_DATA_23_const_net_32             = 4'h0;
assign OE_DATA_24_const_net_32             = 4'h0;
assign OE_DATA_25_const_net_32             = 4'h0;
assign OE_DATA_26_const_net_32             = 4'h0;
assign OE_DATA_27_const_net_32             = 4'h0;
assign OE_DATA_28_const_net_32             = 4'h0;
assign OE_DATA_29_const_net_32             = 4'h0;
assign OE_DATA_30_const_net_32             = 4'h0;
assign OE_DATA_31_const_net_32             = 4'h0;
assign OE_DATA_32_const_net_32             = 4'h0;
assign OE_DATA_33_const_net_32             = 4'h0;
assign OE_DATA_34_const_net_32             = 4'h0;
assign OE_DATA_35_const_net_32             = 4'h0;
assign OE_DATA_36_const_net_32             = 4'h0;
assign OE_DATA_37_const_net_32             = 4'h0;
assign OE_DATA_38_const_net_32             = 4'h0;
assign OE_DATA_39_const_net_32             = 4'h0;
assign OE_DATA_40_const_net_32             = 4'h0;
assign OE_DATA_41_const_net_32             = 4'h0;
assign OE_DATA_42_const_net_32             = 4'h0;
assign OE_DATA_43_const_net_32             = 4'h0;
assign OE_DATA_44_const_net_32             = 4'h0;
assign OE_DATA_45_const_net_32             = 4'h0;
assign OE_DATA_46_const_net_32             = 4'h0;
assign OE_DATA_47_const_net_32             = 4'h0;
assign OE_DATA_48_const_net_32             = 4'h0;
assign OE_DATA_49_const_net_32             = 4'h0;
assign OE_DATA_50_const_net_32             = 4'h0;
assign OE_DATA_51_const_net_32             = 4'h0;
assign OE_DATA_52_const_net_32             = 4'h0;
assign OE_DATA_53_const_net_32             = 4'h0;
assign OE_DATA_54_const_net_32             = 4'h0;
assign OE_DATA_55_const_net_32             = 4'h0;
assign OE_DATA_56_const_net_32             = 4'h0;
assign OE_DATA_57_const_net_32             = 4'h0;
assign OE_DATA_58_const_net_32             = 4'h0;
assign OE_DATA_59_const_net_32             = 4'h0;
assign OE_DATA_60_const_net_32             = 4'h0;
assign OE_DATA_61_const_net_32             = 4'h0;
assign OE_DATA_62_const_net_32             = 4'h0;
assign OE_DATA_63_const_net_32             = 4'h0;
assign OE_DATA_64_const_net_32             = 4'h0;
assign OE_DATA_65_const_net_32             = 4'h0;
assign OE_DATA_66_const_net_32             = 4'h0;
assign OE_DATA_67_const_net_32             = 4'h0;
assign OE_DATA_68_const_net_32             = 4'h0;
assign OE_DATA_69_const_net_32             = 4'h0;
assign OE_DATA_70_const_net_32             = 4'h0;
assign OE_DATA_71_const_net_32             = 4'h0;
assign OE_DATA_72_const_net_32             = 4'h0;
assign OE_DATA_73_const_net_32             = 4'h0;
assign OE_DATA_74_const_net_32             = 4'h0;
assign OE_DATA_75_const_net_32             = 4'h0;
assign OE_DATA_76_const_net_32             = 4'h0;
assign OE_DATA_77_const_net_32             = 4'h0;
assign OE_DATA_78_const_net_32             = 4'h0;
assign OE_DATA_79_const_net_32             = 4'h0;
assign OE_DATA_80_const_net_32             = 4'h0;
assign OE_DATA_81_const_net_32             = 4'h0;
assign OE_DATA_82_const_net_32             = 4'h0;
assign OE_DATA_83_const_net_32             = 4'h0;
assign OE_DATA_84_const_net_32             = 4'h0;
assign OE_DATA_85_const_net_32             = 4'h0;
assign OE_DATA_86_const_net_32             = 4'h0;
assign OE_DATA_87_const_net_32             = 4'h0;
assign OE_DATA_88_const_net_32             = 4'h0;
assign OE_DATA_89_const_net_32             = 4'h0;
assign OE_DATA_90_const_net_32             = 4'h0;
assign OE_DATA_91_const_net_32             = 4'h0;
assign OE_DATA_92_const_net_32             = 4'h0;
assign OE_DATA_93_const_net_32             = 4'h0;
assign OE_DATA_94_const_net_32             = 4'h0;
assign OE_DATA_95_const_net_32             = 4'h0;
assign OE_DATA_96_const_net_32             = 4'h0;
assign OE_DATA_97_const_net_32             = 4'h0;
assign OE_DATA_98_const_net_32             = 4'h0;
assign OE_DATA_99_const_net_32             = 4'h0;
assign OE_DATA_100_const_net_32            = 4'h0;
assign OE_DATA_101_const_net_32            = 4'h0;
assign OE_DATA_102_const_net_32            = 4'h0;
assign OE_DATA_103_const_net_32            = 4'h0;
assign OE_DATA_104_const_net_32            = 4'h0;
assign OE_DATA_105_const_net_32            = 4'h0;
assign OE_DATA_106_const_net_32            = 4'h0;
assign OE_DATA_107_const_net_32            = 4'h0;
assign OE_DATA_108_const_net_32            = 4'h0;
assign OE_DATA_109_const_net_32            = 4'h0;
assign OE_DATA_110_const_net_32            = 4'h0;
assign OE_DATA_111_const_net_32            = 4'h0;
assign OE_DATA_112_const_net_32            = 4'h0;
assign OE_DATA_113_const_net_32            = 4'h0;
assign OE_DATA_114_const_net_32            = 4'h0;
assign OE_DATA_115_const_net_32            = 4'h0;
assign OE_DATA_116_const_net_32            = 4'h0;
assign OE_DATA_117_const_net_32            = 4'h0;
assign OE_DATA_118_const_net_32            = 4'h0;
assign OE_DATA_119_const_net_32            = 4'h0;
assign OE_DATA_120_const_net_32            = 4'h0;
assign OE_DATA_121_const_net_32            = 4'h0;
assign OE_DATA_122_const_net_32            = 4'h0;
assign OE_DATA_123_const_net_32            = 4'h0;
assign OE_DATA_124_const_net_32            = 4'h0;
assign OE_DATA_125_const_net_32            = 4'h0;
assign OE_DATA_126_const_net_32            = 4'h0;
assign OE_DATA_127_const_net_32            = 4'h0;
assign RX_DQS_90_const_net_21              = 2'h0;
assign FIFO_WR_PTR_const_net_22            = 3'h0;
assign FIFO_RD_PTR_const_net_22            = 3'h0;
assign EYE_MONITOR_LANE_WIDTH_const_net_25 = 3'h0;
assign TX_DATA_1_const_net_26              = 2'h0;
assign TX_DATA_2_const_net_28              = 2'h0;
assign TX_DATA_3_const_net_28              = 2'h0;
assign TX_DATA_4_const_net_28              = 2'h0;
assign TX_DATA_5_const_net_28              = 2'h0;
assign TX_DATA_6_const_net_28              = 2'h0;
assign TX_DATA_7_const_net_28              = 2'h0;
assign TX_DATA_8_const_net_32              = 2'h0;
assign TX_DATA_9_const_net_32              = 2'h0;
assign TX_DATA_10_const_net_32             = 2'h0;
assign TX_DATA_11_const_net_32             = 2'h0;
assign TX_DATA_12_const_net_33             = 2'h0;
assign TX_DATA_13_const_net_33             = 2'h0;
assign TX_DATA_14_const_net_33             = 2'h0;
assign TX_DATA_15_const_net_33             = 2'h0;
assign TX_DATA_16_const_net_33             = 2'h0;
assign TX_DATA_17_const_net_33             = 2'h0;
assign TX_DATA_18_const_net_33             = 2'h0;
assign TX_DATA_19_const_net_33             = 2'h0;
assign TX_DATA_20_const_net_33             = 2'h0;
assign TX_DATA_21_const_net_33             = 2'h0;
assign TX_DATA_22_const_net_33             = 2'h0;
assign TX_DATA_23_const_net_33             = 2'h0;
assign TX_DATA_24_const_net_33             = 2'h0;
assign TX_DATA_25_const_net_33             = 2'h0;
assign TX_DATA_26_const_net_33             = 2'h0;
assign TX_DATA_27_const_net_33             = 2'h0;
assign TX_DATA_28_const_net_33             = 2'h0;
assign TX_DATA_29_const_net_33             = 2'h0;
assign TX_DATA_30_const_net_33             = 2'h0;
assign TX_DATA_31_const_net_33             = 2'h0;
assign TX_DATA_32_const_net_33             = 2'h0;
assign TX_DATA_33_const_net_33             = 2'h0;
assign TX_DATA_34_const_net_33             = 2'h0;
assign TX_DATA_35_const_net_33             = 2'h0;
assign TX_DATA_36_const_net_33             = 2'h0;
assign TX_DATA_37_const_net_33             = 2'h0;
assign TX_DATA_38_const_net_33             = 2'h0;
assign TX_DATA_39_const_net_33             = 2'h0;
assign TX_DATA_40_const_net_33             = 2'h0;
assign TX_DATA_41_const_net_33             = 2'h0;
assign TX_DATA_42_const_net_33             = 2'h0;
assign TX_DATA_43_const_net_33             = 2'h0;
assign TX_DATA_44_const_net_33             = 2'h0;
assign TX_DATA_45_const_net_33             = 2'h0;
assign TX_DATA_46_const_net_33             = 2'h0;
assign TX_DATA_47_const_net_33             = 2'h0;
assign TX_DATA_48_const_net_33             = 2'h0;
assign TX_DATA_49_const_net_33             = 2'h0;
assign TX_DATA_50_const_net_33             = 2'h0;
assign TX_DATA_51_const_net_33             = 2'h0;
assign TX_DATA_52_const_net_33             = 2'h0;
assign TX_DATA_53_const_net_33             = 2'h0;
assign TX_DATA_54_const_net_33             = 2'h0;
assign TX_DATA_55_const_net_33             = 2'h0;
assign TX_DATA_56_const_net_33             = 2'h0;
assign TX_DATA_57_const_net_33             = 2'h0;
assign TX_DATA_58_const_net_33             = 2'h0;
assign TX_DATA_59_const_net_33             = 2'h0;
assign TX_DATA_60_const_net_33             = 2'h0;
assign TX_DATA_61_const_net_33             = 2'h0;
assign TX_DATA_62_const_net_33             = 2'h0;
assign TX_DATA_63_const_net_33             = 2'h0;
assign TX_DATA_64_const_net_33             = 2'h0;
assign TX_DATA_65_const_net_33             = 2'h0;
assign TX_DATA_66_const_net_33             = 2'h0;
assign TX_DATA_67_const_net_33             = 2'h0;
assign TX_DATA_68_const_net_33             = 2'h0;
assign TX_DATA_69_const_net_33             = 2'h0;
assign TX_DATA_70_const_net_33             = 2'h0;
assign TX_DATA_71_const_net_33             = 2'h0;
assign TX_DATA_72_const_net_33             = 2'h0;
assign TX_DATA_73_const_net_33             = 2'h0;
assign TX_DATA_74_const_net_33             = 2'h0;
assign TX_DATA_75_const_net_33             = 2'h0;
assign TX_DATA_76_const_net_33             = 2'h0;
assign TX_DATA_77_const_net_33             = 2'h0;
assign TX_DATA_78_const_net_33             = 2'h0;
assign TX_DATA_79_const_net_33             = 2'h0;
assign TX_DATA_80_const_net_33             = 2'h0;
assign TX_DATA_81_const_net_33             = 2'h0;
assign TX_DATA_82_const_net_33             = 2'h0;
assign TX_DATA_83_const_net_33             = 2'h0;
assign TX_DATA_84_const_net_33             = 2'h0;
assign TX_DATA_85_const_net_33             = 2'h0;
assign TX_DATA_86_const_net_33             = 2'h0;
assign TX_DATA_87_const_net_33             = 2'h0;
assign TX_DATA_88_const_net_33             = 2'h0;
assign TX_DATA_89_const_net_33             = 2'h0;
assign TX_DATA_90_const_net_33             = 2'h0;
assign TX_DATA_91_const_net_33             = 2'h0;
assign TX_DATA_92_const_net_33             = 2'h0;
assign TX_DATA_93_const_net_33             = 2'h0;
assign TX_DATA_94_const_net_33             = 2'h0;
assign TX_DATA_95_const_net_33             = 2'h0;
assign TX_DATA_96_const_net_33             = 2'h0;
assign TX_DATA_97_const_net_33             = 2'h0;
assign TX_DATA_98_const_net_33             = 2'h0;
assign TX_DATA_99_const_net_33             = 2'h0;
assign TX_DATA_100_const_net_33            = 2'h0;
assign TX_DATA_101_const_net_33            = 2'h0;
assign TX_DATA_102_const_net_33            = 2'h0;
assign TX_DATA_103_const_net_33            = 2'h0;
assign TX_DATA_104_const_net_33            = 2'h0;
assign TX_DATA_105_const_net_33            = 2'h0;
assign TX_DATA_106_const_net_33            = 2'h0;
assign TX_DATA_107_const_net_33            = 2'h0;
assign TX_DATA_108_const_net_33            = 2'h0;
assign TX_DATA_109_const_net_33            = 2'h0;
assign TX_DATA_110_const_net_33            = 2'h0;
assign TX_DATA_111_const_net_33            = 2'h0;
assign TX_DATA_112_const_net_33            = 2'h0;
assign TX_DATA_113_const_net_33            = 2'h0;
assign TX_DATA_114_const_net_33            = 2'h0;
assign TX_DATA_115_const_net_33            = 2'h0;
assign TX_DATA_116_const_net_33            = 2'h0;
assign TX_DATA_117_const_net_33            = 2'h0;
assign TX_DATA_118_const_net_33            = 2'h0;
assign TX_DATA_119_const_net_33            = 2'h0;
assign TX_DATA_120_const_net_33            = 2'h0;
assign TX_DATA_121_const_net_33            = 2'h0;
assign TX_DATA_122_const_net_33            = 2'h0;
assign TX_DATA_123_const_net_33            = 2'h0;
assign TX_DATA_124_const_net_33            = 2'h0;
assign TX_DATA_125_const_net_33            = 2'h0;
assign TX_DATA_126_const_net_33            = 2'h0;
assign TX_DATA_127_const_net_33            = 2'h0;
assign OE_DATA_1_const_net_29              = 2'h0;
assign OE_DATA_2_const_net_29              = 2'h0;
assign OE_DATA_3_const_net_29              = 2'h0;
assign OE_DATA_4_const_net_29              = 2'h0;
assign OE_DATA_5_const_net_29              = 2'h0;
assign OE_DATA_6_const_net_29              = 2'h0;
assign OE_DATA_7_const_net_29              = 2'h0;
assign OE_DATA_8_const_net_33              = 2'h0;
assign OE_DATA_9_const_net_33              = 2'h0;
assign OE_DATA_10_const_net_33             = 2'h0;
assign OE_DATA_11_const_net_33             = 2'h0;
assign OE_DATA_12_const_net_33             = 2'h0;
assign OE_DATA_13_const_net_33             = 2'h0;
assign OE_DATA_14_const_net_33             = 2'h0;
assign OE_DATA_15_const_net_33             = 2'h0;
assign OE_DATA_16_const_net_33             = 2'h0;
assign OE_DATA_17_const_net_33             = 2'h0;
assign OE_DATA_18_const_net_33             = 2'h0;
assign OE_DATA_19_const_net_33             = 2'h0;
assign OE_DATA_20_const_net_33             = 2'h0;
assign OE_DATA_21_const_net_33             = 2'h0;
assign OE_DATA_22_const_net_33             = 2'h0;
assign OE_DATA_23_const_net_33             = 2'h0;
assign OE_DATA_24_const_net_33             = 2'h0;
assign OE_DATA_25_const_net_33             = 2'h0;
assign OE_DATA_26_const_net_33             = 2'h0;
assign OE_DATA_27_const_net_33             = 2'h0;
assign OE_DATA_28_const_net_33             = 2'h0;
assign OE_DATA_29_const_net_33             = 2'h0;
assign OE_DATA_30_const_net_33             = 2'h0;
assign OE_DATA_31_const_net_33             = 2'h0;
assign OE_DATA_32_const_net_33             = 2'h0;
assign OE_DATA_33_const_net_33             = 2'h0;
assign OE_DATA_34_const_net_33             = 2'h0;
assign OE_DATA_35_const_net_33             = 2'h0;
assign OE_DATA_36_const_net_33             = 2'h0;
assign OE_DATA_37_const_net_33             = 2'h0;
assign OE_DATA_38_const_net_33             = 2'h0;
assign OE_DATA_39_const_net_33             = 2'h0;
assign OE_DATA_40_const_net_33             = 2'h0;
assign OE_DATA_41_const_net_33             = 2'h0;
assign OE_DATA_42_const_net_33             = 2'h0;
assign OE_DATA_43_const_net_33             = 2'h0;
assign OE_DATA_44_const_net_33             = 2'h0;
assign OE_DATA_45_const_net_33             = 2'h0;
assign OE_DATA_46_const_net_33             = 2'h0;
assign OE_DATA_47_const_net_33             = 2'h0;
assign OE_DATA_48_const_net_33             = 2'h0;
assign OE_DATA_49_const_net_33             = 2'h0;
assign OE_DATA_50_const_net_33             = 2'h0;
assign OE_DATA_51_const_net_33             = 2'h0;
assign OE_DATA_52_const_net_33             = 2'h0;
assign OE_DATA_53_const_net_33             = 2'h0;
assign OE_DATA_54_const_net_33             = 2'h0;
assign OE_DATA_55_const_net_33             = 2'h0;
assign OE_DATA_56_const_net_33             = 2'h0;
assign OE_DATA_57_const_net_33             = 2'h0;
assign OE_DATA_58_const_net_33             = 2'h0;
assign OE_DATA_59_const_net_33             = 2'h0;
assign OE_DATA_60_const_net_33             = 2'h0;
assign OE_DATA_61_const_net_33             = 2'h0;
assign OE_DATA_62_const_net_33             = 2'h0;
assign OE_DATA_63_const_net_33             = 2'h0;
assign OE_DATA_64_const_net_33             = 2'h0;
assign OE_DATA_65_const_net_33             = 2'h0;
assign OE_DATA_66_const_net_33             = 2'h0;
assign OE_DATA_67_const_net_33             = 2'h0;
assign OE_DATA_68_const_net_33             = 2'h0;
assign OE_DATA_69_const_net_33             = 2'h0;
assign OE_DATA_70_const_net_33             = 2'h0;
assign OE_DATA_71_const_net_33             = 2'h0;
assign OE_DATA_72_const_net_33             = 2'h0;
assign OE_DATA_73_const_net_33             = 2'h0;
assign OE_DATA_74_const_net_33             = 2'h0;
assign OE_DATA_75_const_net_33             = 2'h0;
assign OE_DATA_76_const_net_33             = 2'h0;
assign OE_DATA_77_const_net_33             = 2'h0;
assign OE_DATA_78_const_net_33             = 2'h0;
assign OE_DATA_79_const_net_33             = 2'h0;
assign OE_DATA_80_const_net_33             = 2'h0;
assign OE_DATA_81_const_net_33             = 2'h0;
assign OE_DATA_82_const_net_33             = 2'h0;
assign OE_DATA_83_const_net_33             = 2'h0;
assign OE_DATA_84_const_net_33             = 2'h0;
assign OE_DATA_85_const_net_33             = 2'h0;
assign OE_DATA_86_const_net_33             = 2'h0;
assign OE_DATA_87_const_net_33             = 2'h0;
assign OE_DATA_88_const_net_33             = 2'h0;
assign OE_DATA_89_const_net_33             = 2'h0;
assign OE_DATA_90_const_net_33             = 2'h0;
assign OE_DATA_91_const_net_33             = 2'h0;
assign OE_DATA_92_const_net_33             = 2'h0;
assign OE_DATA_93_const_net_33             = 2'h0;
assign OE_DATA_94_const_net_33             = 2'h0;
assign OE_DATA_95_const_net_33             = 2'h0;
assign OE_DATA_96_const_net_33             = 2'h0;
assign OE_DATA_97_const_net_33             = 2'h0;
assign OE_DATA_98_const_net_33             = 2'h0;
assign OE_DATA_99_const_net_33             = 2'h0;
assign OE_DATA_100_const_net_33            = 2'h0;
assign OE_DATA_101_const_net_33            = 2'h0;
assign OE_DATA_102_const_net_33            = 2'h0;
assign OE_DATA_103_const_net_33            = 2'h0;
assign OE_DATA_104_const_net_33            = 2'h0;
assign OE_DATA_105_const_net_33            = 2'h0;
assign OE_DATA_106_const_net_33            = 2'h0;
assign OE_DATA_107_const_net_33            = 2'h0;
assign OE_DATA_108_const_net_33            = 2'h0;
assign OE_DATA_109_const_net_33            = 2'h0;
assign OE_DATA_110_const_net_33            = 2'h0;
assign OE_DATA_111_const_net_33            = 2'h0;
assign OE_DATA_112_const_net_33            = 2'h0;
assign OE_DATA_113_const_net_33            = 2'h0;
assign OE_DATA_114_const_net_33            = 2'h0;
assign OE_DATA_115_const_net_33            = 2'h0;
assign OE_DATA_116_const_net_33            = 2'h0;
assign OE_DATA_117_const_net_33            = 2'h0;
assign OE_DATA_118_const_net_33            = 2'h0;
assign OE_DATA_119_const_net_33            = 2'h0;
assign OE_DATA_120_const_net_33            = 2'h0;
assign OE_DATA_121_const_net_33            = 2'h0;
assign OE_DATA_122_const_net_33            = 2'h0;
assign OE_DATA_123_const_net_33            = 2'h0;
assign OE_DATA_124_const_net_33            = 2'h0;
assign OE_DATA_125_const_net_33            = 2'h0;
assign OE_DATA_126_const_net_33            = 2'h0;
assign OE_DATA_127_const_net_33            = 2'h0;
assign RX_DQS_90_const_net_22              = 2'h0;
assign EYE_MONITOR_LANE_WIDTH_const_net_26 = 3'h0;
assign TX_DATA_1_const_net_27              = 8'h00;
assign TX_DATA_2_const_net_29              = 8'h00;
assign TX_DATA_3_const_net_29              = 8'h00;
assign TX_DATA_4_const_net_29              = 8'h00;
assign TX_DATA_5_const_net_29              = 8'h00;
assign TX_DATA_6_const_net_29              = 8'h00;
assign TX_DATA_7_const_net_29              = 8'h00;
assign TX_DATA_8_const_net_33              = 8'h00;
assign TX_DATA_9_const_net_33              = 8'h00;
assign TX_DATA_10_const_net_33             = 8'h00;
assign TX_DATA_11_const_net_33             = 8'h00;
assign TX_DATA_12_const_net_34             = 8'h00;
assign TX_DATA_13_const_net_34             = 8'h00;
assign TX_DATA_14_const_net_34             = 8'h00;
assign TX_DATA_15_const_net_34             = 8'h00;
assign TX_DATA_16_const_net_34             = 8'h00;
assign TX_DATA_17_const_net_34             = 8'h00;
assign TX_DATA_18_const_net_34             = 8'h00;
assign TX_DATA_19_const_net_34             = 8'h00;
assign TX_DATA_20_const_net_34             = 8'h00;
assign TX_DATA_21_const_net_34             = 8'h00;
assign TX_DATA_22_const_net_34             = 8'h00;
assign TX_DATA_23_const_net_34             = 8'h00;
assign TX_DATA_24_const_net_34             = 8'h00;
assign TX_DATA_25_const_net_34             = 8'h00;
assign TX_DATA_26_const_net_34             = 8'h00;
assign TX_DATA_27_const_net_34             = 8'h00;
assign TX_DATA_28_const_net_34             = 8'h00;
assign TX_DATA_29_const_net_34             = 8'h00;
assign TX_DATA_30_const_net_34             = 8'h00;
assign TX_DATA_31_const_net_34             = 8'h00;
assign TX_DATA_32_const_net_34             = 8'h00;
assign TX_DATA_33_const_net_34             = 8'h00;
assign TX_DATA_34_const_net_34             = 8'h00;
assign TX_DATA_35_const_net_34             = 8'h00;
assign TX_DATA_36_const_net_34             = 8'h00;
assign TX_DATA_37_const_net_34             = 8'h00;
assign TX_DATA_38_const_net_34             = 8'h00;
assign TX_DATA_39_const_net_34             = 8'h00;
assign TX_DATA_40_const_net_34             = 8'h00;
assign TX_DATA_41_const_net_34             = 8'h00;
assign TX_DATA_42_const_net_34             = 8'h00;
assign TX_DATA_43_const_net_34             = 8'h00;
assign TX_DATA_44_const_net_34             = 8'h00;
assign TX_DATA_45_const_net_34             = 8'h00;
assign TX_DATA_46_const_net_34             = 8'h00;
assign TX_DATA_47_const_net_34             = 8'h00;
assign TX_DATA_48_const_net_34             = 8'h00;
assign TX_DATA_49_const_net_34             = 8'h00;
assign TX_DATA_50_const_net_34             = 8'h00;
assign TX_DATA_51_const_net_34             = 8'h00;
assign TX_DATA_52_const_net_34             = 8'h00;
assign TX_DATA_53_const_net_34             = 8'h00;
assign TX_DATA_54_const_net_34             = 8'h00;
assign TX_DATA_55_const_net_34             = 8'h00;
assign TX_DATA_56_const_net_34             = 8'h00;
assign TX_DATA_57_const_net_34             = 8'h00;
assign TX_DATA_58_const_net_34             = 8'h00;
assign TX_DATA_59_const_net_34             = 8'h00;
assign TX_DATA_60_const_net_34             = 8'h00;
assign TX_DATA_61_const_net_34             = 8'h00;
assign TX_DATA_62_const_net_34             = 8'h00;
assign TX_DATA_63_const_net_34             = 8'h00;
assign TX_DATA_64_const_net_34             = 8'h00;
assign TX_DATA_65_const_net_34             = 8'h00;
assign TX_DATA_66_const_net_34             = 8'h00;
assign TX_DATA_67_const_net_34             = 8'h00;
assign TX_DATA_68_const_net_34             = 8'h00;
assign TX_DATA_69_const_net_34             = 8'h00;
assign TX_DATA_70_const_net_34             = 8'h00;
assign TX_DATA_71_const_net_34             = 8'h00;
assign TX_DATA_72_const_net_34             = 8'h00;
assign TX_DATA_73_const_net_34             = 8'h00;
assign TX_DATA_74_const_net_34             = 8'h00;
assign TX_DATA_75_const_net_34             = 8'h00;
assign TX_DATA_76_const_net_34             = 8'h00;
assign TX_DATA_77_const_net_34             = 8'h00;
assign TX_DATA_78_const_net_34             = 8'h00;
assign TX_DATA_79_const_net_34             = 8'h00;
assign TX_DATA_80_const_net_34             = 8'h00;
assign TX_DATA_81_const_net_34             = 8'h00;
assign TX_DATA_82_const_net_34             = 8'h00;
assign TX_DATA_83_const_net_34             = 8'h00;
assign TX_DATA_84_const_net_34             = 8'h00;
assign TX_DATA_85_const_net_34             = 8'h00;
assign TX_DATA_86_const_net_34             = 8'h00;
assign TX_DATA_87_const_net_34             = 8'h00;
assign TX_DATA_88_const_net_34             = 8'h00;
assign TX_DATA_89_const_net_34             = 8'h00;
assign TX_DATA_90_const_net_34             = 8'h00;
assign TX_DATA_91_const_net_34             = 8'h00;
assign TX_DATA_92_const_net_34             = 8'h00;
assign TX_DATA_93_const_net_34             = 8'h00;
assign TX_DATA_94_const_net_34             = 8'h00;
assign TX_DATA_95_const_net_34             = 8'h00;
assign TX_DATA_96_const_net_34             = 8'h00;
assign TX_DATA_97_const_net_34             = 8'h00;
assign TX_DATA_98_const_net_34             = 8'h00;
assign TX_DATA_99_const_net_34             = 8'h00;
assign TX_DATA_100_const_net_34            = 8'h00;
assign TX_DATA_101_const_net_34            = 8'h00;
assign TX_DATA_102_const_net_34            = 8'h00;
assign TX_DATA_103_const_net_34            = 8'h00;
assign TX_DATA_104_const_net_34            = 8'h00;
assign TX_DATA_105_const_net_34            = 8'h00;
assign TX_DATA_106_const_net_34            = 8'h00;
assign TX_DATA_107_const_net_34            = 8'h00;
assign TX_DATA_108_const_net_34            = 8'h00;
assign TX_DATA_109_const_net_34            = 8'h00;
assign TX_DATA_110_const_net_34            = 8'h00;
assign TX_DATA_111_const_net_34            = 8'h00;
assign TX_DATA_112_const_net_34            = 8'h00;
assign TX_DATA_113_const_net_34            = 8'h00;
assign TX_DATA_114_const_net_34            = 8'h00;
assign TX_DATA_115_const_net_34            = 8'h00;
assign TX_DATA_116_const_net_34            = 8'h00;
assign TX_DATA_117_const_net_34            = 8'h00;
assign TX_DATA_118_const_net_34            = 8'h00;
assign TX_DATA_119_const_net_34            = 8'h00;
assign TX_DATA_120_const_net_34            = 8'h00;
assign TX_DATA_121_const_net_34            = 8'h00;
assign TX_DATA_122_const_net_34            = 8'h00;
assign TX_DATA_123_const_net_34            = 8'h00;
assign TX_DATA_124_const_net_34            = 8'h00;
assign TX_DATA_125_const_net_34            = 8'h00;
assign TX_DATA_126_const_net_34            = 8'h00;
assign TX_DATA_127_const_net_34            = 8'h00;
assign OE_DATA_1_const_net_30              = 4'h0;
assign OE_DATA_2_const_net_30              = 4'h0;
assign OE_DATA_3_const_net_30              = 4'h0;
assign OE_DATA_4_const_net_30              = 4'h0;
assign OE_DATA_5_const_net_30              = 4'h0;
assign OE_DATA_6_const_net_30              = 4'h0;
assign OE_DATA_7_const_net_30              = 4'h0;
assign OE_DATA_8_const_net_34              = 4'h0;
assign OE_DATA_9_const_net_34              = 4'h0;
assign OE_DATA_10_const_net_34             = 4'h0;
assign OE_DATA_11_const_net_34             = 4'h0;
assign OE_DATA_12_const_net_34             = 4'h0;
assign OE_DATA_13_const_net_34             = 4'h0;
assign OE_DATA_14_const_net_34             = 4'h0;
assign OE_DATA_15_const_net_34             = 4'h0;
assign OE_DATA_16_const_net_34             = 4'h0;
assign OE_DATA_17_const_net_34             = 4'h0;
assign OE_DATA_18_const_net_34             = 4'h0;
assign OE_DATA_19_const_net_34             = 4'h0;
assign OE_DATA_20_const_net_34             = 4'h0;
assign OE_DATA_21_const_net_34             = 4'h0;
assign OE_DATA_22_const_net_34             = 4'h0;
assign OE_DATA_23_const_net_34             = 4'h0;
assign OE_DATA_24_const_net_34             = 4'h0;
assign OE_DATA_25_const_net_34             = 4'h0;
assign OE_DATA_26_const_net_34             = 4'h0;
assign OE_DATA_27_const_net_34             = 4'h0;
assign OE_DATA_28_const_net_34             = 4'h0;
assign OE_DATA_29_const_net_34             = 4'h0;
assign OE_DATA_30_const_net_34             = 4'h0;
assign OE_DATA_31_const_net_34             = 4'h0;
assign OE_DATA_32_const_net_34             = 4'h0;
assign OE_DATA_33_const_net_34             = 4'h0;
assign OE_DATA_34_const_net_34             = 4'h0;
assign OE_DATA_35_const_net_34             = 4'h0;
assign OE_DATA_36_const_net_34             = 4'h0;
assign OE_DATA_37_const_net_34             = 4'h0;
assign OE_DATA_38_const_net_34             = 4'h0;
assign OE_DATA_39_const_net_34             = 4'h0;
assign OE_DATA_40_const_net_34             = 4'h0;
assign OE_DATA_41_const_net_34             = 4'h0;
assign OE_DATA_42_const_net_34             = 4'h0;
assign OE_DATA_43_const_net_34             = 4'h0;
assign OE_DATA_44_const_net_34             = 4'h0;
assign OE_DATA_45_const_net_34             = 4'h0;
assign OE_DATA_46_const_net_34             = 4'h0;
assign OE_DATA_47_const_net_34             = 4'h0;
assign OE_DATA_48_const_net_34             = 4'h0;
assign OE_DATA_49_const_net_34             = 4'h0;
assign OE_DATA_50_const_net_34             = 4'h0;
assign OE_DATA_51_const_net_34             = 4'h0;
assign OE_DATA_52_const_net_34             = 4'h0;
assign OE_DATA_53_const_net_34             = 4'h0;
assign OE_DATA_54_const_net_34             = 4'h0;
assign OE_DATA_55_const_net_34             = 4'h0;
assign OE_DATA_56_const_net_34             = 4'h0;
assign OE_DATA_57_const_net_34             = 4'h0;
assign OE_DATA_58_const_net_34             = 4'h0;
assign OE_DATA_59_const_net_34             = 4'h0;
assign OE_DATA_60_const_net_34             = 4'h0;
assign OE_DATA_61_const_net_34             = 4'h0;
assign OE_DATA_62_const_net_34             = 4'h0;
assign OE_DATA_63_const_net_34             = 4'h0;
assign OE_DATA_64_const_net_34             = 4'h0;
assign OE_DATA_65_const_net_34             = 4'h0;
assign OE_DATA_66_const_net_34             = 4'h0;
assign OE_DATA_67_const_net_34             = 4'h0;
assign OE_DATA_68_const_net_34             = 4'h0;
assign OE_DATA_69_const_net_34             = 4'h0;
assign OE_DATA_70_const_net_34             = 4'h0;
assign OE_DATA_71_const_net_34             = 4'h0;
assign OE_DATA_72_const_net_34             = 4'h0;
assign OE_DATA_73_const_net_34             = 4'h0;
assign OE_DATA_74_const_net_34             = 4'h0;
assign OE_DATA_75_const_net_34             = 4'h0;
assign OE_DATA_76_const_net_34             = 4'h0;
assign OE_DATA_77_const_net_34             = 4'h0;
assign OE_DATA_78_const_net_34             = 4'h0;
assign OE_DATA_79_const_net_34             = 4'h0;
assign OE_DATA_80_const_net_34             = 4'h0;
assign OE_DATA_81_const_net_34             = 4'h0;
assign OE_DATA_82_const_net_34             = 4'h0;
assign OE_DATA_83_const_net_34             = 4'h0;
assign OE_DATA_84_const_net_34             = 4'h0;
assign OE_DATA_85_const_net_34             = 4'h0;
assign OE_DATA_86_const_net_34             = 4'h0;
assign OE_DATA_87_const_net_34             = 4'h0;
assign OE_DATA_88_const_net_34             = 4'h0;
assign OE_DATA_89_const_net_34             = 4'h0;
assign OE_DATA_90_const_net_34             = 4'h0;
assign OE_DATA_91_const_net_34             = 4'h0;
assign OE_DATA_92_const_net_34             = 4'h0;
assign OE_DATA_93_const_net_34             = 4'h0;
assign OE_DATA_94_const_net_34             = 4'h0;
assign OE_DATA_95_const_net_34             = 4'h0;
assign OE_DATA_96_const_net_34             = 4'h0;
assign OE_DATA_97_const_net_34             = 4'h0;
assign OE_DATA_98_const_net_34             = 4'h0;
assign OE_DATA_99_const_net_34             = 4'h0;
assign OE_DATA_100_const_net_34            = 4'h0;
assign OE_DATA_101_const_net_34            = 4'h0;
assign OE_DATA_102_const_net_34            = 4'h0;
assign OE_DATA_103_const_net_34            = 4'h0;
assign OE_DATA_104_const_net_34            = 4'h0;
assign OE_DATA_105_const_net_34            = 4'h0;
assign OE_DATA_106_const_net_34            = 4'h0;
assign OE_DATA_107_const_net_34            = 4'h0;
assign OE_DATA_108_const_net_34            = 4'h0;
assign OE_DATA_109_const_net_34            = 4'h0;
assign OE_DATA_110_const_net_34            = 4'h0;
assign OE_DATA_111_const_net_34            = 4'h0;
assign OE_DATA_112_const_net_34            = 4'h0;
assign OE_DATA_113_const_net_34            = 4'h0;
assign OE_DATA_114_const_net_34            = 4'h0;
assign OE_DATA_115_const_net_34            = 4'h0;
assign OE_DATA_116_const_net_34            = 4'h0;
assign OE_DATA_117_const_net_34            = 4'h0;
assign OE_DATA_118_const_net_34            = 4'h0;
assign OE_DATA_119_const_net_34            = 4'h0;
assign OE_DATA_120_const_net_34            = 4'h0;
assign OE_DATA_121_const_net_34            = 4'h0;
assign OE_DATA_122_const_net_34            = 4'h0;
assign OE_DATA_123_const_net_34            = 4'h0;
assign OE_DATA_124_const_net_34            = 4'h0;
assign OE_DATA_125_const_net_34            = 4'h0;
assign OE_DATA_126_const_net_34            = 4'h0;
assign OE_DATA_127_const_net_34            = 4'h0;
assign READ_CLK_SEL_const_net_0            = 3'h0;
assign EYE_MONITOR_WIDTH_IN_const_net_4    = 3'h0;
assign CDR_CLK_A_SEL_const_net_0           = 8'h00;
assign CDR_CLK_B_SEL_const_net_4           = 11'h000;
//--------------------------------------------------------------------
// Inversions
//--------------------------------------------------------------------
assign SYNC_SYS_RST_N_net_1 = ~ SYNC_SYS_RST_N_OUT_PRE_INV0_0;
//--------------------------------------------------------------------
// TieOff assignments
//--------------------------------------------------------------------
assign DFI_CALVL_RESP[1:0]           = 2'h0;
assign DFI_CALVL_TRAIN_DONE          = 1'b1;
assign DFI_CTRLUPD_ACK               = 1'b0;
assign DFI_PHYUPD_REQ                = 1'b0;
assign DFI_PHYUPD_TYPE[1:0]          = 2'h0;
//--------------------------------------------------------------------
// Top level output port assignments
//--------------------------------------------------------------------
assign CODE_UPDATE_net_1             = CODE_UPDATE_net_0;
assign CODE_UPDATE                   = CODE_UPDATE_net_1;
assign LOADPHS_B_net_1[0]            = LOADPHS_B_net_0[0];
assign LOADPHS_B[0:0]                = LOADPHS_B_net_1[0];
assign VCO_PHSEL_BCLK_SEL_net_1[0]   = VCO_PHSEL_BCLK_SEL_net_0[0];
assign VCO_PHSEL_BCLK_SEL[0:0]       = VCO_PHSEL_BCLK_SEL_net_1[0];
assign VCO_PHSEL_BCLK90_SEL_net_1[0] = VCO_PHSEL_BCLK90_SEL_net_0[0];
assign VCO_PHSEL_BCLK90_SEL[0:0]     = VCO_PHSEL_BCLK90_SEL_net_1[0];
assign VCO_PHSEL_REFCLK_SEL_net_1    = VCO_PHSEL_REFCLK_SEL_net_0;
assign VCO_PHSEL_REFCLK_SEL          = VCO_PHSEL_REFCLK_SEL_net_1;
assign VCO_PHSEL_ROTATE_net_1[0]     = VCO_PHSEL_ROTATE_net_0[0];
assign VCO_PHSEL_ROTATE[0:0]         = VCO_PHSEL_ROTATE_net_1[0];
assign DFI_RDDATA_W0_net_1           = DFI_RDDATA_W0_net_0;
assign DFI_RDDATA_W0[63:0]           = DFI_RDDATA_W0_net_1;
assign DFI_RDDATA_VALID_W0_net_1[0]  = DFI_RDDATA_VALID_W0_net_0;
assign DFI_RDDATA_VALID_W0[0:0]      = DFI_RDDATA_VALID_W0_net_1[0];
assign DFI_RDDATA_VALID_W0_net_2[1]  = DFI_RDDATA_VALID_W0_net_0;
assign DFI_RDDATA_VALID_W0[1:1]      = DFI_RDDATA_VALID_W0_net_2[1];
assign DFI_RDDATA_VALID_W0_net_3[2]  = DFI_RDDATA_VALID_W0_net_0;
assign DFI_RDDATA_VALID_W0[2:2]      = DFI_RDDATA_VALID_W0_net_3[2];
assign DFI_RDDATA_VALID_W0_net_4[3]  = DFI_RDDATA_VALID_W0_net_0;
assign DFI_RDDATA_VALID_W0[3:3]      = DFI_RDDATA_VALID_W0_net_4[3];
assign DFI_RDDATA_W1_net_1           = DFI_RDDATA_W1_net_0;
assign DFI_RDDATA_W1[63:0]           = DFI_RDDATA_W1_net_1;
assign DFI_RDDATA_VALID_W1_net_1[0]  = DFI_RDDATA_VALID_W1_net_0;
assign DFI_RDDATA_VALID_W1[0:0]      = DFI_RDDATA_VALID_W1_net_1[0];
assign DFI_RDDATA_VALID_W1_net_2[1]  = DFI_RDDATA_VALID_W1_net_0;
assign DFI_RDDATA_VALID_W1[1:1]      = DFI_RDDATA_VALID_W1_net_2[1];
assign DFI_RDDATA_VALID_W1_net_3[2]  = DFI_RDDATA_VALID_W1_net_0;
assign DFI_RDDATA_VALID_W1[2:2]      = DFI_RDDATA_VALID_W1_net_3[2];
assign DFI_RDDATA_VALID_W1_net_4[3]  = DFI_RDDATA_VALID_W1_net_0;
assign DFI_RDDATA_VALID_W1[3:3]      = DFI_RDDATA_VALID_W1_net_4[3];
assign DFI_RDDATA_W2_net_1           = DFI_RDDATA_W2_net_0;
assign DFI_RDDATA_W2[63:0]           = DFI_RDDATA_W2_net_1;
assign DFI_RDDATA_VALID_W2_net_1[0]  = DFI_RDDATA_VALID_W2_net_0;
assign DFI_RDDATA_VALID_W2[0:0]      = DFI_RDDATA_VALID_W2_net_1[0];
assign DFI_RDDATA_VALID_W2_net_2[1]  = DFI_RDDATA_VALID_W2_net_0;
assign DFI_RDDATA_VALID_W2[1:1]      = DFI_RDDATA_VALID_W2_net_2[1];
assign DFI_RDDATA_VALID_W2_net_3[2]  = DFI_RDDATA_VALID_W2_net_0;
assign DFI_RDDATA_VALID_W2[2:2]      = DFI_RDDATA_VALID_W2_net_3[2];
assign DFI_RDDATA_VALID_W2_net_4[3]  = DFI_RDDATA_VALID_W2_net_0;
assign DFI_RDDATA_VALID_W2[3:3]      = DFI_RDDATA_VALID_W2_net_4[3];
assign DFI_RDDATA_W3_net_1           = DFI_RDDATA_W3_net_0;
assign DFI_RDDATA_W3[63:0]           = DFI_RDDATA_W3_net_1;
assign DFI_RDDATA_VALID_W3_net_1[0]  = DFI_RDDATA_VALID_W3_net_0;
assign DFI_RDDATA_VALID_W3[0:0]      = DFI_RDDATA_VALID_W3_net_1[0];
assign DFI_RDDATA_VALID_W3_net_2[1]  = DFI_RDDATA_VALID_W3_net_0;
assign DFI_RDDATA_VALID_W3[1:1]      = DFI_RDDATA_VALID_W3_net_2[1];
assign DFI_RDDATA_VALID_W3_net_3[2]  = DFI_RDDATA_VALID_W3_net_0;
assign DFI_RDDATA_VALID_W3[2:2]      = DFI_RDDATA_VALID_W3_net_3[2];
assign DFI_RDDATA_VALID_W3_net_4[3]  = DFI_RDDATA_VALID_W3_net_0;
assign DFI_RDDATA_VALID_W3[3:3]      = DFI_RDDATA_VALID_W3_net_4[3];
assign DFI_RDLVL_RESP_net_1          = DFI_RDLVL_RESP_net_0;
assign DFI_RDLVL_RESP[3:0]           = DFI_RDLVL_RESP_net_1;
assign DFI_WRLVL_RESP_net_1          = DFI_WRLVL_RESP_net_0;
assign DFI_WRLVL_RESP[3:0]           = DFI_WRLVL_RESP_net_1;
assign DFI_INIT_COMPLETE_net_1       = DFI_INIT_COMPLETE_net_0;
assign DFI_INIT_COMPLETE             = DFI_INIT_COMPLETE_net_1;
assign DFI_TRAINING_COMPLETE_net_1   = DFI_TRAINING_COMPLETE_net_0;
assign DFI_TRAINING_COMPLETE         = DFI_TRAINING_COMPLETE_net_1;
assign DM_N_net_1[0]                 = DM_N_net_0[0];
assign DM_N[0:0]                     = DM_N_net_1[0];
assign DM_N_0_net_0[1]               = DM_N_0[0];
assign DM_N[1:1]                     = DM_N_0_net_0[1];
assign DM_N_1_net_0[2]               = DM_N_1[0];
assign DM_N[2:2]                     = DM_N_1_net_0[2];
assign DM_N_2_net_0[3]               = DM_N_2[0];
assign DM_N[3:3]                     = DM_N_2_net_0[3];
assign CKE_net_1                     = CKE_net_0[0];
assign CKE                           = CKE_net_1;
assign CS_N_net_1                    = CS_N_net_0[0];
assign CS_N                          = CS_N_net_1;
assign ODT_net_1                     = ODT_net_0[0];
assign ODT                           = ODT_net_1;
assign RAS_N_net_1                   = RAS_N_net_0[0];
assign RAS_N                         = RAS_N_net_1;
assign CAS_N_net_1                   = CAS_N_net_0[0];
assign CAS_N                         = CAS_N_net_1;
assign WE_N_net_1                    = WE_N_net_0[0];
assign WE_N                          = WE_N_net_1;
assign ACT_N_net_1                   = ACT_N_net_0[0];
assign ACT_N                         = ACT_N_net_1;
assign BG_net_1                      = BG_net_0;
assign BG[1:0]                       = BG_net_1;
assign BA_net_1                      = BA_net_0;
assign BA[1:0]                       = BA_net_1;
assign RESET_N_net_1                 = RESET_N_net_0[0];
assign RESET_N                       = RESET_N_net_1;
assign A_net_1[0]                    = A_net_0[0];
assign A[0:0]                        = A_net_1[0];
assign A_9_net_0[10]                 = A_9[10];
assign A[10:10]                      = A_9_net_0[10];
assign A_10_net_0[11]                = A_10[11];
assign A[11:11]                      = A_10_net_0[11];
assign A_11_net_0[12]                = A_11;
assign A[12:12]                      = A_11_net_0[12];
assign A_12_net_0[13]                = A_12[0];
assign A[13:13]                      = A_12_net_0[13];
assign A_0_net_0[1]                  = A_0[1];
assign A[1:1]                        = A_0_net_0[1];
assign A_1_net_0[2]                  = A_1[2];
assign A[2:2]                        = A_1_net_0[2];
assign A_2_net_0[3]                  = A_2[3];
assign A[3:3]                        = A_2_net_0[3];
assign A_3_net_0[4]                  = A_3[4];
assign A[4:4]                        = A_3_net_0[4];
assign A_4_net_0[5]                  = A_4[5];
assign A[5:5]                        = A_4_net_0[5];
assign A_5_net_0[6]                  = A_5[6];
assign A[6:6]                        = A_5_net_0[6];
assign A_6_net_0[7]                  = A_6[7];
assign A[7:7]                        = A_6_net_0[7];
assign A_7_net_0[8]                  = A_7[8];
assign A[8:8]                        = A_7_net_0[8];
assign A_8_net_0[9]                  = A_8[9];
assign A[9:9]                        = A_8_net_0[9];
assign CK0_net_1                     = CK0_net_0;
assign CK0                           = CK0_net_1;
assign CK0_N_net_1                   = CK0_N_net_0;
assign CK0_N                         = CK0_N_net_1;
assign SHIELD0_net_1                 = SHIELD0_net_0;
assign SHIELD0                       = SHIELD0_net_1;
assign SHIELD1_net_1                 = SHIELD1_net_0;
assign SHIELD1                       = SHIELD1_net_1;
assign SHIELD2_net_1                 = SHIELD2_net_0;
assign SHIELD2                       = SHIELD2_net_1;
assign SHIELD3_net_1                 = SHIELD3_net_0;
assign SHIELD3                       = SHIELD3_net_1;
assign APB_DEBUG_PRDATA_net_0        = APB_DEBUG_PRDATA;
assign PRDATA[7:0]                   = APB_DEBUG_PRDATA_net_0;
assign APB_DEBUG_PREADY_net_0        = APB_DEBUG_PREADY;
assign PREADY                        = APB_DEBUG_PREADY_net_0;
assign CAL_INIT_MR_W_REQ_net_1       = CAL_INIT_MR_W_REQ_net_0;
assign CAL_INIT_MR_W_REQ             = CAL_INIT_MR_W_REQ_net_1;
assign CAL_INIT_MR_ADDR_net_1        = CAL_INIT_MR_ADDR_net_0;
assign CAL_INIT_MR_ADDR[7:0]         = CAL_INIT_MR_ADDR_net_1;
assign CAL_INIT_MR_WR_DATA_net_1     = CAL_INIT_MR_WR_DATA_net_0;
assign CAL_INIT_MR_WR_DATA[17:0]     = CAL_INIT_MR_WR_DATA_net_1;
assign CAL_INIT_MR_WR_MASK_net_1     = CAL_INIT_MR_WR_MASK_net_0;
assign CAL_INIT_MR_WR_MASK[17:0]     = CAL_INIT_MR_WR_MASK_net_1;
assign CAL_INIT_CS_net_1             = CAL_INIT_CS_net_0;
assign CAL_INIT_CS[1:0]              = CAL_INIT_CS_net_1;
assign CTRLR_READY_OUT_net_1         = CTRLR_READY_OUT_net_0;
assign CTRLR_READY_OUT               = CTRLR_READY_OUT_net_1;
assign ITER_COUNT_net_1              = ITER_COUNT_net_0;
assign ITER_COUNT[3:0]               = ITER_COUNT_net_1;
assign CAL_L_R_REQ_net_1             = CAL_L_R_REQ_net_0;
assign CAL_L_R_REQ                   = CAL_L_R_REQ_net_1;
assign CAL_L_W_REQ_net_1             = CAL_L_W_REQ_net_0;
assign CAL_L_W_REQ                   = CAL_L_W_REQ_net_1;
assign CAL_L_DATAIN_net_1            = CAL_L_DATAIN_net_0;
assign CAL_L_DATAIN[255:0]           = CAL_L_DATAIN_net_1;
assign CAL_L_DM_IN_net_1             = CAL_L_DM_IN_net_0;
assign CAL_L_DM_IN[31:0]             = CAL_L_DM_IN_net_1;
assign CAL_SELECT_net_1              = CAL_SELECT_net_0;
assign CAL_SELECT                    = CAL_SELECT_net_1;
assign SYNC_SYS_RST_N_OUT_PRE_INV0_0 = SYNC_SYS_RST_N_net_0;
assign SYNC_SYS_RST_N                = SYNC_SYS_RST_N_net_1;
//--------------------------------------------------------------------
// Slices assignments
//--------------------------------------------------------------------
assign A_net_0[0]                                          = PAD_O_net_0[0:0];
assign A_0[1]                                              = PAD_O_net_0[1:1];
assign A_1[2]                                              = PAD_O_net_0[2:2];
assign A_2[3]                                              = PAD_O_net_0[3:3];
assign A_3[4]                                              = PAD_O_net_0[4:4];
assign A_4[5]                                              = PAD_O_net_0[5:5];
assign A_5[6]                                              = PAD_O_net_0[6:6];
assign A_6[7]                                              = PAD_O_net_0[7:7];
assign A_7[8]                                              = PAD_O_net_0[8:8];
assign A_8[9]                                              = PAD_O_net_0[9:9];
assign A_9[10]                                             = PAD_O_net_0[10:10];
assign A_10[11]                                            = PAD_O_net_0[11:11];
assign DFI_ADDRESS_P0_slice_0[0]                           = DFI_ADDRESS_P0[0:0];
assign DFI_ADDRESS_P0_slice_1[1]                           = DFI_ADDRESS_P0[1:1];
assign DFI_ADDRESS_P0_slice_2[2]                           = DFI_ADDRESS_P0[2:2];
assign DFI_ADDRESS_P0_slice_3[3]                           = DFI_ADDRESS_P0[3:3];
assign DFI_ADDRESS_P0_slice_4[4]                           = DFI_ADDRESS_P0[4:4];
assign DFI_ADDRESS_P0_slice_5[5]                           = DFI_ADDRESS_P0[5:5];
assign DFI_ADDRESS_P0_slice_6[6]                           = DFI_ADDRESS_P0[6:6];
assign DFI_ADDRESS_P0_slice_7[7]                           = DFI_ADDRESS_P0[7:7];
assign DFI_ADDRESS_P0_slice_8[8]                           = DFI_ADDRESS_P0[8:8];
assign DFI_ADDRESS_P0_slice_9[9]                           = DFI_ADDRESS_P0[9:9];
assign DFI_ADDRESS_P0_slice_10[10]                         = DFI_ADDRESS_P0[10:10];
assign DFI_ADDRESS_P0_slice_11[11]                         = DFI_ADDRESS_P0[11:11];
assign DFI_ADDRESS_P0_slice_12[12]                         = DFI_ADDRESS_P0[12:12];
assign DFI_ADDRESS_P0_slice_13[13]                         = DFI_ADDRESS_P0[13:13];
assign DFI_ADDRESS_P1_slice_0[0]                           = DFI_ADDRESS_P1[0:0];
assign DFI_ADDRESS_P1_slice_1[1]                           = DFI_ADDRESS_P1[1:1];
assign DFI_ADDRESS_P1_slice_2[2]                           = DFI_ADDRESS_P1[2:2];
assign DFI_ADDRESS_P1_slice_3[3]                           = DFI_ADDRESS_P1[3:3];
assign DFI_ADDRESS_P1_slice_4[4]                           = DFI_ADDRESS_P1[4:4];
assign DFI_ADDRESS_P1_slice_5[5]                           = DFI_ADDRESS_P1[5:5];
assign DFI_ADDRESS_P1_slice_6[6]                           = DFI_ADDRESS_P1[6:6];
assign DFI_ADDRESS_P1_slice_7[7]                           = DFI_ADDRESS_P1[7:7];
assign DFI_ADDRESS_P1_slice_8[8]                           = DFI_ADDRESS_P1[8:8];
assign DFI_ADDRESS_P1_slice_9[9]                           = DFI_ADDRESS_P1[9:9];
assign DFI_ADDRESS_P1_slice_10[10]                         = DFI_ADDRESS_P1[10:10];
assign DFI_ADDRESS_P1_slice_11[11]                         = DFI_ADDRESS_P1[11:11];
assign DFI_ADDRESS_P1_slice_12[12]                         = DFI_ADDRESS_P1[12:12];
assign DFI_ADDRESS_P1_slice_13[13]                         = DFI_ADDRESS_P1[13:13];
assign DFI_ADDRESS_P2_slice_0[0]                           = DFI_ADDRESS_P2[0:0];
assign DFI_ADDRESS_P2_slice_1[1]                           = DFI_ADDRESS_P2[1:1];
assign DFI_ADDRESS_P2_slice_2[2]                           = DFI_ADDRESS_P2[2:2];
assign DFI_ADDRESS_P2_slice_3[3]                           = DFI_ADDRESS_P2[3:3];
assign DFI_ADDRESS_P2_slice_4[4]                           = DFI_ADDRESS_P2[4:4];
assign DFI_ADDRESS_P2_slice_5[5]                           = DFI_ADDRESS_P2[5:5];
assign DFI_ADDRESS_P2_slice_6[6]                           = DFI_ADDRESS_P2[6:6];
assign DFI_ADDRESS_P2_slice_7[7]                           = DFI_ADDRESS_P2[7:7];
assign DFI_ADDRESS_P2_slice_8[8]                           = DFI_ADDRESS_P2[8:8];
assign DFI_ADDRESS_P2_slice_9[9]                           = DFI_ADDRESS_P2[9:9];
assign DFI_ADDRESS_P2_slice_10[10]                         = DFI_ADDRESS_P2[10:10];
assign DFI_ADDRESS_P2_slice_11[11]                         = DFI_ADDRESS_P2[11:11];
assign DFI_ADDRESS_P2_slice_12[12]                         = DFI_ADDRESS_P2[12:12];
assign DFI_ADDRESS_P2_slice_13[13]                         = DFI_ADDRESS_P2[13:13];
assign DFI_ADDRESS_P3_slice_0[0]                           = DFI_ADDRESS_P3[0:0];
assign DFI_ADDRESS_P3_slice_1[1]                           = DFI_ADDRESS_P3[1:1];
assign DFI_ADDRESS_P3_slice_2[2]                           = DFI_ADDRESS_P3[2:2];
assign DFI_ADDRESS_P3_slice_3[3]                           = DFI_ADDRESS_P3[3:3];
assign DFI_ADDRESS_P3_slice_4[4]                           = DFI_ADDRESS_P3[4:4];
assign DFI_ADDRESS_P3_slice_5[5]                           = DFI_ADDRESS_P3[5:5];
assign DFI_ADDRESS_P3_slice_6[6]                           = DFI_ADDRESS_P3[6:6];
assign DFI_ADDRESS_P3_slice_7[7]                           = DFI_ADDRESS_P3[7:7];
assign DFI_ADDRESS_P3_slice_8[8]                           = DFI_ADDRESS_P3[8:8];
assign DFI_ADDRESS_P3_slice_9[9]                           = DFI_ADDRESS_P3[9:9];
assign DFI_ADDRESS_P3_slice_10[10]                         = DFI_ADDRESS_P3[10:10];
assign DFI_ADDRESS_P3_slice_11[11]                         = DFI_ADDRESS_P3[11:11];
assign DFI_ADDRESS_P3_slice_12[12]                         = DFI_ADDRESS_P3[12:12];
assign DFI_ADDRESS_P3_slice_13[13]                         = DFI_ADDRESS_P3[13:13];
assign DFI_BANK_P0_slice_0[0]                              = DFI_BANK_P0[0:0];
assign DFI_BANK_P0_slice_1[1]                              = DFI_BANK_P0[1:1];
assign DFI_BANK_P1_slice_0[0]                              = DFI_BANK_P1[0:0];
assign DFI_BANK_P1_slice_1[1]                              = DFI_BANK_P1[1:1];
assign DFI_BANK_P2_slice_0[0]                              = DFI_BANK_P2[0:0];
assign DFI_BANK_P2_slice_1[1]                              = DFI_BANK_P2[1:1];
assign DFI_BANK_P3_slice_0[0]                              = DFI_BANK_P3[0:0];
assign DFI_BANK_P3_slice_1[1]                              = DFI_BANK_P3[1:1];
assign DFI_BG_P0_slice_0[0]                                = DFI_BG_P0[0:0];
assign DFI_BG_P0_slice_1[1]                                = DFI_BG_P0[1:1];
assign DFI_BG_P1_slice_0[0]                                = DFI_BG_P1[0:0];
assign DFI_BG_P1_slice_1[1]                                = DFI_BG_P1[1:1];
assign DFI_BG_P2_slice_0[0]                                = DFI_BG_P2[0:0];
assign DFI_BG_P2_slice_1[1]                                = DFI_BG_P2[1:1];
assign DFI_BG_P3_slice_0[0]                                = DFI_BG_P3[0:0];
assign DFI_BG_P3_slice_1[1]                                = DFI_BG_P3[1:1];
assign DFI_RDDATA_EN_P0_slice_0[0]                         = DFI_RDDATA_EN_P0[0:0];
assign DFI_RDDATA_EN_P1_slice_0[0]                         = DFI_RDDATA_EN_P1[0:0];
assign DFI_RDDATA_EN_P2_slice_0[0]                         = DFI_RDDATA_EN_P2[0:0];
assign DFI_RDDATA_EN_P3_slice_0[0]                         = DFI_RDDATA_EN_P3[0:0];
assign DFI_WRDATA_EN_P0_slice_0[0]                         = DFI_WRDATA_EN_P0[0:0];
assign DFI_WRDATA_EN_P1_slice_0[0]                         = DFI_WRDATA_EN_P1[0:0];
assign DFI_WRDATA_EN_P2_slice_0[0]                         = DFI_WRDATA_EN_P2[0:0];
assign DFI_WRDATA_EN_P3_slice_0[0]                         = DFI_WRDATA_EN_P3[0:0];
assign DFI_WRDATA_MASK_P0_slice_0[0]                       = DFI_WRDATA_MASK_P0[0:0];
assign DFI_WRDATA_MASK_P0_slice_1[4]                       = DFI_WRDATA_MASK_P0[4:4];
assign DFI_WRDATA_MASK_P0_slice_2[1]                       = DFI_WRDATA_MASK_P0[1:1];
assign DFI_WRDATA_MASK_P0_slice_3[5]                       = DFI_WRDATA_MASK_P0[5:5];
assign DFI_WRDATA_MASK_P0_slice_4[2]                       = DFI_WRDATA_MASK_P0[2:2];
assign DFI_WRDATA_MASK_P0_slice_5[6]                       = DFI_WRDATA_MASK_P0[6:6];
assign DFI_WRDATA_MASK_P0_slice_6[3]                       = DFI_WRDATA_MASK_P0[3:3];
assign DFI_WRDATA_MASK_P0_slice_7[7]                       = DFI_WRDATA_MASK_P0[7:7];
assign DFI_WRDATA_MASK_P1_slice_0[0]                       = DFI_WRDATA_MASK_P1[0:0];
assign DFI_WRDATA_MASK_P1_slice_1[4]                       = DFI_WRDATA_MASK_P1[4:4];
assign DFI_WRDATA_MASK_P1_slice_2[1]                       = DFI_WRDATA_MASK_P1[1:1];
assign DFI_WRDATA_MASK_P1_slice_3[5]                       = DFI_WRDATA_MASK_P1[5:5];
assign DFI_WRDATA_MASK_P1_slice_4[2]                       = DFI_WRDATA_MASK_P1[2:2];
assign DFI_WRDATA_MASK_P1_slice_5[6]                       = DFI_WRDATA_MASK_P1[6:6];
assign DFI_WRDATA_MASK_P1_slice_6[3]                       = DFI_WRDATA_MASK_P1[3:3];
assign DFI_WRDATA_MASK_P1_slice_7[7]                       = DFI_WRDATA_MASK_P1[7:7];
assign DFI_WRDATA_MASK_P2_slice_0[0]                       = DFI_WRDATA_MASK_P2[0:0];
assign DFI_WRDATA_MASK_P2_slice_1[4]                       = DFI_WRDATA_MASK_P2[4:4];
assign DFI_WRDATA_MASK_P2_slice_2[1]                       = DFI_WRDATA_MASK_P2[1:1];
assign DFI_WRDATA_MASK_P2_slice_3[5]                       = DFI_WRDATA_MASK_P2[5:5];
assign DFI_WRDATA_MASK_P2_slice_4[2]                       = DFI_WRDATA_MASK_P2[2:2];
assign DFI_WRDATA_MASK_P2_slice_5[6]                       = DFI_WRDATA_MASK_P2[6:6];
assign DFI_WRDATA_MASK_P2_slice_6[3]                       = DFI_WRDATA_MASK_P2[3:3];
assign DFI_WRDATA_MASK_P2_slice_7[7]                       = DFI_WRDATA_MASK_P2[7:7];
assign DFI_WRDATA_MASK_P3_slice_0[0]                       = DFI_WRDATA_MASK_P3[0:0];
assign DFI_WRDATA_MASK_P3_slice_1[4]                       = DFI_WRDATA_MASK_P3[4:4];
assign DFI_WRDATA_MASK_P3_slice_2[1]                       = DFI_WRDATA_MASK_P3[1:1];
assign DFI_WRDATA_MASK_P3_slice_3[5]                       = DFI_WRDATA_MASK_P3[5:5];
assign DFI_WRDATA_MASK_P3_slice_4[2]                       = DFI_WRDATA_MASK_P3[2:2];
assign DFI_WRDATA_MASK_P3_slice_5[6]                       = DFI_WRDATA_MASK_P3[6:6];
assign DFI_WRDATA_MASK_P3_slice_6[3]                       = DFI_WRDATA_MASK_P3[3:3];
assign DFI_WRDATA_MASK_P3_slice_7[7]                       = DFI_WRDATA_MASK_P3[7:7];
assign DFI_WRDATA_P0_slice_0[0]                            = DFI_WRDATA_P0[0:0];
assign DFI_WRDATA_P0_slice_1[32]                           = DFI_WRDATA_P0[32:32];
assign DFI_WRDATA_P0_slice_2[1]                            = DFI_WRDATA_P0[1:1];
assign DFI_WRDATA_P0_slice_3[33]                           = DFI_WRDATA_P0[33:33];
assign DFI_WRDATA_P0_slice_4[2]                            = DFI_WRDATA_P0[2:2];
assign DFI_WRDATA_P0_slice_5[34]                           = DFI_WRDATA_P0[34:34];
assign DFI_WRDATA_P0_slice_6[3]                            = DFI_WRDATA_P0[3:3];
assign DFI_WRDATA_P0_slice_7[35]                           = DFI_WRDATA_P0[35:35];
assign DFI_WRDATA_P0_slice_8[4]                            = DFI_WRDATA_P0[4:4];
assign DFI_WRDATA_P0_slice_9[36]                           = DFI_WRDATA_P0[36:36];
assign DFI_WRDATA_P0_slice_10[5]                           = DFI_WRDATA_P0[5:5];
assign DFI_WRDATA_P0_slice_11[37]                          = DFI_WRDATA_P0[37:37];
assign DFI_WRDATA_P0_slice_12[6]                           = DFI_WRDATA_P0[6:6];
assign DFI_WRDATA_P0_slice_13[38]                          = DFI_WRDATA_P0[38:38];
assign DFI_WRDATA_P0_slice_14[7]                           = DFI_WRDATA_P0[7:7];
assign DFI_WRDATA_P0_slice_15[39]                          = DFI_WRDATA_P0[39:39];
assign DFI_WRDATA_P0_slice_16[8]                           = DFI_WRDATA_P0[8:8];
assign DFI_WRDATA_P0_slice_17[40]                          = DFI_WRDATA_P0[40:40];
assign DFI_WRDATA_P0_slice_18[9]                           = DFI_WRDATA_P0[9:9];
assign DFI_WRDATA_P0_slice_19[41]                          = DFI_WRDATA_P0[41:41];
assign DFI_WRDATA_P0_slice_20[10]                          = DFI_WRDATA_P0[10:10];
assign DFI_WRDATA_P0_slice_21[42]                          = DFI_WRDATA_P0[42:42];
assign DFI_WRDATA_P0_slice_22[11]                          = DFI_WRDATA_P0[11:11];
assign DFI_WRDATA_P0_slice_23[43]                          = DFI_WRDATA_P0[43:43];
assign DFI_WRDATA_P0_slice_24[12]                          = DFI_WRDATA_P0[12:12];
assign DFI_WRDATA_P0_slice_25[44]                          = DFI_WRDATA_P0[44:44];
assign DFI_WRDATA_P0_slice_26[13]                          = DFI_WRDATA_P0[13:13];
assign DFI_WRDATA_P0_slice_27[45]                          = DFI_WRDATA_P0[45:45];
assign DFI_WRDATA_P0_slice_28[14]                          = DFI_WRDATA_P0[14:14];
assign DFI_WRDATA_P0_slice_29[46]                          = DFI_WRDATA_P0[46:46];
assign DFI_WRDATA_P0_slice_30[15]                          = DFI_WRDATA_P0[15:15];
assign DFI_WRDATA_P0_slice_31[47]                          = DFI_WRDATA_P0[47:47];
assign DFI_WRDATA_P0_slice_32[16]                          = DFI_WRDATA_P0[16:16];
assign DFI_WRDATA_P0_slice_33[48]                          = DFI_WRDATA_P0[48:48];
assign DFI_WRDATA_P0_slice_34[17]                          = DFI_WRDATA_P0[17:17];
assign DFI_WRDATA_P0_slice_35[49]                          = DFI_WRDATA_P0[49:49];
assign DFI_WRDATA_P0_slice_36[18]                          = DFI_WRDATA_P0[18:18];
assign DFI_WRDATA_P0_slice_37[50]                          = DFI_WRDATA_P0[50:50];
assign DFI_WRDATA_P0_slice_38[19]                          = DFI_WRDATA_P0[19:19];
assign DFI_WRDATA_P0_slice_39[51]                          = DFI_WRDATA_P0[51:51];
assign DFI_WRDATA_P0_slice_40[20]                          = DFI_WRDATA_P0[20:20];
assign DFI_WRDATA_P0_slice_41[52]                          = DFI_WRDATA_P0[52:52];
assign DFI_WRDATA_P0_slice_42[21]                          = DFI_WRDATA_P0[21:21];
assign DFI_WRDATA_P0_slice_43[53]                          = DFI_WRDATA_P0[53:53];
assign DFI_WRDATA_P0_slice_44[22]                          = DFI_WRDATA_P0[22:22];
assign DFI_WRDATA_P0_slice_45[54]                          = DFI_WRDATA_P0[54:54];
assign DFI_WRDATA_P0_slice_46[23]                          = DFI_WRDATA_P0[23:23];
assign DFI_WRDATA_P0_slice_47[55]                          = DFI_WRDATA_P0[55:55];
assign DFI_WRDATA_P0_slice_48[24]                          = DFI_WRDATA_P0[24:24];
assign DFI_WRDATA_P0_slice_49[56]                          = DFI_WRDATA_P0[56:56];
assign DFI_WRDATA_P0_slice_50[25]                          = DFI_WRDATA_P0[25:25];
assign DFI_WRDATA_P0_slice_51[57]                          = DFI_WRDATA_P0[57:57];
assign DFI_WRDATA_P0_slice_52[26]                          = DFI_WRDATA_P0[26:26];
assign DFI_WRDATA_P0_slice_53[58]                          = DFI_WRDATA_P0[58:58];
assign DFI_WRDATA_P0_slice_54[27]                          = DFI_WRDATA_P0[27:27];
assign DFI_WRDATA_P0_slice_55[59]                          = DFI_WRDATA_P0[59:59];
assign DFI_WRDATA_P0_slice_56[28]                          = DFI_WRDATA_P0[28:28];
assign DFI_WRDATA_P0_slice_57[60]                          = DFI_WRDATA_P0[60:60];
assign DFI_WRDATA_P0_slice_58[29]                          = DFI_WRDATA_P0[29:29];
assign DFI_WRDATA_P0_slice_59[61]                          = DFI_WRDATA_P0[61:61];
assign DFI_WRDATA_P0_slice_60[30]                          = DFI_WRDATA_P0[30:30];
assign DFI_WRDATA_P0_slice_61[62]                          = DFI_WRDATA_P0[62:62];
assign DFI_WRDATA_P0_slice_62[31]                          = DFI_WRDATA_P0[31:31];
assign DFI_WRDATA_P0_slice_63[63]                          = DFI_WRDATA_P0[63:63];
assign DFI_WRDATA_P1_slice_0[0]                            = DFI_WRDATA_P1[0:0];
assign DFI_WRDATA_P1_slice_1[32]                           = DFI_WRDATA_P1[32:32];
assign DFI_WRDATA_P1_slice_2[1]                            = DFI_WRDATA_P1[1:1];
assign DFI_WRDATA_P1_slice_3[33]                           = DFI_WRDATA_P1[33:33];
assign DFI_WRDATA_P1_slice_4[2]                            = DFI_WRDATA_P1[2:2];
assign DFI_WRDATA_P1_slice_5[34]                           = DFI_WRDATA_P1[34:34];
assign DFI_WRDATA_P1_slice_6[3]                            = DFI_WRDATA_P1[3:3];
assign DFI_WRDATA_P1_slice_7[35]                           = DFI_WRDATA_P1[35:35];
assign DFI_WRDATA_P1_slice_8[4]                            = DFI_WRDATA_P1[4:4];
assign DFI_WRDATA_P1_slice_9[36]                           = DFI_WRDATA_P1[36:36];
assign DFI_WRDATA_P1_slice_10[5]                           = DFI_WRDATA_P1[5:5];
assign DFI_WRDATA_P1_slice_11[37]                          = DFI_WRDATA_P1[37:37];
assign DFI_WRDATA_P1_slice_12[6]                           = DFI_WRDATA_P1[6:6];
assign DFI_WRDATA_P1_slice_13[38]                          = DFI_WRDATA_P1[38:38];
assign DFI_WRDATA_P1_slice_14[7]                           = DFI_WRDATA_P1[7:7];
assign DFI_WRDATA_P1_slice_15[39]                          = DFI_WRDATA_P1[39:39];
assign DFI_WRDATA_P1_slice_16[8]                           = DFI_WRDATA_P1[8:8];
assign DFI_WRDATA_P1_slice_17[40]                          = DFI_WRDATA_P1[40:40];
assign DFI_WRDATA_P1_slice_18[9]                           = DFI_WRDATA_P1[9:9];
assign DFI_WRDATA_P1_slice_19[41]                          = DFI_WRDATA_P1[41:41];
assign DFI_WRDATA_P1_slice_20[10]                          = DFI_WRDATA_P1[10:10];
assign DFI_WRDATA_P1_slice_21[42]                          = DFI_WRDATA_P1[42:42];
assign DFI_WRDATA_P1_slice_22[11]                          = DFI_WRDATA_P1[11:11];
assign DFI_WRDATA_P1_slice_23[43]                          = DFI_WRDATA_P1[43:43];
assign DFI_WRDATA_P1_slice_24[12]                          = DFI_WRDATA_P1[12:12];
assign DFI_WRDATA_P1_slice_25[44]                          = DFI_WRDATA_P1[44:44];
assign DFI_WRDATA_P1_slice_26[13]                          = DFI_WRDATA_P1[13:13];
assign DFI_WRDATA_P1_slice_27[45]                          = DFI_WRDATA_P1[45:45];
assign DFI_WRDATA_P1_slice_28[14]                          = DFI_WRDATA_P1[14:14];
assign DFI_WRDATA_P1_slice_29[46]                          = DFI_WRDATA_P1[46:46];
assign DFI_WRDATA_P1_slice_30[15]                          = DFI_WRDATA_P1[15:15];
assign DFI_WRDATA_P1_slice_31[47]                          = DFI_WRDATA_P1[47:47];
assign DFI_WRDATA_P1_slice_32[16]                          = DFI_WRDATA_P1[16:16];
assign DFI_WRDATA_P1_slice_33[48]                          = DFI_WRDATA_P1[48:48];
assign DFI_WRDATA_P1_slice_34[17]                          = DFI_WRDATA_P1[17:17];
assign DFI_WRDATA_P1_slice_35[49]                          = DFI_WRDATA_P1[49:49];
assign DFI_WRDATA_P1_slice_36[18]                          = DFI_WRDATA_P1[18:18];
assign DFI_WRDATA_P1_slice_37[50]                          = DFI_WRDATA_P1[50:50];
assign DFI_WRDATA_P1_slice_38[19]                          = DFI_WRDATA_P1[19:19];
assign DFI_WRDATA_P1_slice_39[51]                          = DFI_WRDATA_P1[51:51];
assign DFI_WRDATA_P1_slice_40[20]                          = DFI_WRDATA_P1[20:20];
assign DFI_WRDATA_P1_slice_41[52]                          = DFI_WRDATA_P1[52:52];
assign DFI_WRDATA_P1_slice_42[21]                          = DFI_WRDATA_P1[21:21];
assign DFI_WRDATA_P1_slice_43[53]                          = DFI_WRDATA_P1[53:53];
assign DFI_WRDATA_P1_slice_44[22]                          = DFI_WRDATA_P1[22:22];
assign DFI_WRDATA_P1_slice_45[54]                          = DFI_WRDATA_P1[54:54];
assign DFI_WRDATA_P1_slice_46[23]                          = DFI_WRDATA_P1[23:23];
assign DFI_WRDATA_P1_slice_47[55]                          = DFI_WRDATA_P1[55:55];
assign DFI_WRDATA_P1_slice_48[24]                          = DFI_WRDATA_P1[24:24];
assign DFI_WRDATA_P1_slice_49[56]                          = DFI_WRDATA_P1[56:56];
assign DFI_WRDATA_P1_slice_50[25]                          = DFI_WRDATA_P1[25:25];
assign DFI_WRDATA_P1_slice_51[57]                          = DFI_WRDATA_P1[57:57];
assign DFI_WRDATA_P1_slice_52[26]                          = DFI_WRDATA_P1[26:26];
assign DFI_WRDATA_P1_slice_53[58]                          = DFI_WRDATA_P1[58:58];
assign DFI_WRDATA_P1_slice_54[27]                          = DFI_WRDATA_P1[27:27];
assign DFI_WRDATA_P1_slice_55[59]                          = DFI_WRDATA_P1[59:59];
assign DFI_WRDATA_P1_slice_56[28]                          = DFI_WRDATA_P1[28:28];
assign DFI_WRDATA_P1_slice_57[60]                          = DFI_WRDATA_P1[60:60];
assign DFI_WRDATA_P1_slice_58[29]                          = DFI_WRDATA_P1[29:29];
assign DFI_WRDATA_P1_slice_59[61]                          = DFI_WRDATA_P1[61:61];
assign DFI_WRDATA_P1_slice_60[30]                          = DFI_WRDATA_P1[30:30];
assign DFI_WRDATA_P1_slice_61[62]                          = DFI_WRDATA_P1[62:62];
assign DFI_WRDATA_P1_slice_62[31]                          = DFI_WRDATA_P1[31:31];
assign DFI_WRDATA_P1_slice_63[63]                          = DFI_WRDATA_P1[63:63];
assign DFI_WRDATA_P2_slice_0[0]                            = DFI_WRDATA_P2[0:0];
assign DFI_WRDATA_P2_slice_1[32]                           = DFI_WRDATA_P2[32:32];
assign DFI_WRDATA_P2_slice_2[1]                            = DFI_WRDATA_P2[1:1];
assign DFI_WRDATA_P2_slice_3[33]                           = DFI_WRDATA_P2[33:33];
assign DFI_WRDATA_P2_slice_4[2]                            = DFI_WRDATA_P2[2:2];
assign DFI_WRDATA_P2_slice_5[34]                           = DFI_WRDATA_P2[34:34];
assign DFI_WRDATA_P2_slice_6[3]                            = DFI_WRDATA_P2[3:3];
assign DFI_WRDATA_P2_slice_7[35]                           = DFI_WRDATA_P2[35:35];
assign DFI_WRDATA_P2_slice_8[4]                            = DFI_WRDATA_P2[4:4];
assign DFI_WRDATA_P2_slice_9[36]                           = DFI_WRDATA_P2[36:36];
assign DFI_WRDATA_P2_slice_10[5]                           = DFI_WRDATA_P2[5:5];
assign DFI_WRDATA_P2_slice_11[37]                          = DFI_WRDATA_P2[37:37];
assign DFI_WRDATA_P2_slice_12[6]                           = DFI_WRDATA_P2[6:6];
assign DFI_WRDATA_P2_slice_13[38]                          = DFI_WRDATA_P2[38:38];
assign DFI_WRDATA_P2_slice_14[7]                           = DFI_WRDATA_P2[7:7];
assign DFI_WRDATA_P2_slice_15[39]                          = DFI_WRDATA_P2[39:39];
assign DFI_WRDATA_P2_slice_16[8]                           = DFI_WRDATA_P2[8:8];
assign DFI_WRDATA_P2_slice_17[40]                          = DFI_WRDATA_P2[40:40];
assign DFI_WRDATA_P2_slice_18[9]                           = DFI_WRDATA_P2[9:9];
assign DFI_WRDATA_P2_slice_19[41]                          = DFI_WRDATA_P2[41:41];
assign DFI_WRDATA_P2_slice_20[10]                          = DFI_WRDATA_P2[10:10];
assign DFI_WRDATA_P2_slice_21[42]                          = DFI_WRDATA_P2[42:42];
assign DFI_WRDATA_P2_slice_22[11]                          = DFI_WRDATA_P2[11:11];
assign DFI_WRDATA_P2_slice_23[43]                          = DFI_WRDATA_P2[43:43];
assign DFI_WRDATA_P2_slice_24[12]                          = DFI_WRDATA_P2[12:12];
assign DFI_WRDATA_P2_slice_25[44]                          = DFI_WRDATA_P2[44:44];
assign DFI_WRDATA_P2_slice_26[13]                          = DFI_WRDATA_P2[13:13];
assign DFI_WRDATA_P2_slice_27[45]                          = DFI_WRDATA_P2[45:45];
assign DFI_WRDATA_P2_slice_28[14]                          = DFI_WRDATA_P2[14:14];
assign DFI_WRDATA_P2_slice_29[46]                          = DFI_WRDATA_P2[46:46];
assign DFI_WRDATA_P2_slice_30[15]                          = DFI_WRDATA_P2[15:15];
assign DFI_WRDATA_P2_slice_31[47]                          = DFI_WRDATA_P2[47:47];
assign DFI_WRDATA_P2_slice_32[16]                          = DFI_WRDATA_P2[16:16];
assign DFI_WRDATA_P2_slice_33[48]                          = DFI_WRDATA_P2[48:48];
assign DFI_WRDATA_P2_slice_34[17]                          = DFI_WRDATA_P2[17:17];
assign DFI_WRDATA_P2_slice_35[49]                          = DFI_WRDATA_P2[49:49];
assign DFI_WRDATA_P2_slice_36[18]                          = DFI_WRDATA_P2[18:18];
assign DFI_WRDATA_P2_slice_37[50]                          = DFI_WRDATA_P2[50:50];
assign DFI_WRDATA_P2_slice_38[19]                          = DFI_WRDATA_P2[19:19];
assign DFI_WRDATA_P2_slice_39[51]                          = DFI_WRDATA_P2[51:51];
assign DFI_WRDATA_P2_slice_40[20]                          = DFI_WRDATA_P2[20:20];
assign DFI_WRDATA_P2_slice_41[52]                          = DFI_WRDATA_P2[52:52];
assign DFI_WRDATA_P2_slice_42[21]                          = DFI_WRDATA_P2[21:21];
assign DFI_WRDATA_P2_slice_43[53]                          = DFI_WRDATA_P2[53:53];
assign DFI_WRDATA_P2_slice_44[22]                          = DFI_WRDATA_P2[22:22];
assign DFI_WRDATA_P2_slice_45[54]                          = DFI_WRDATA_P2[54:54];
assign DFI_WRDATA_P2_slice_46[23]                          = DFI_WRDATA_P2[23:23];
assign DFI_WRDATA_P2_slice_47[55]                          = DFI_WRDATA_P2[55:55];
assign DFI_WRDATA_P2_slice_48[24]                          = DFI_WRDATA_P2[24:24];
assign DFI_WRDATA_P2_slice_49[56]                          = DFI_WRDATA_P2[56:56];
assign DFI_WRDATA_P2_slice_50[25]                          = DFI_WRDATA_P2[25:25];
assign DFI_WRDATA_P2_slice_51[57]                          = DFI_WRDATA_P2[57:57];
assign DFI_WRDATA_P2_slice_52[26]                          = DFI_WRDATA_P2[26:26];
assign DFI_WRDATA_P2_slice_53[58]                          = DFI_WRDATA_P2[58:58];
assign DFI_WRDATA_P2_slice_54[27]                          = DFI_WRDATA_P2[27:27];
assign DFI_WRDATA_P2_slice_55[59]                          = DFI_WRDATA_P2[59:59];
assign DFI_WRDATA_P2_slice_56[28]                          = DFI_WRDATA_P2[28:28];
assign DFI_WRDATA_P2_slice_57[60]                          = DFI_WRDATA_P2[60:60];
assign DFI_WRDATA_P2_slice_58[29]                          = DFI_WRDATA_P2[29:29];
assign DFI_WRDATA_P2_slice_59[61]                          = DFI_WRDATA_P2[61:61];
assign DFI_WRDATA_P2_slice_60[30]                          = DFI_WRDATA_P2[30:30];
assign DFI_WRDATA_P2_slice_61[62]                          = DFI_WRDATA_P2[62:62];
assign DFI_WRDATA_P2_slice_62[31]                          = DFI_WRDATA_P2[31:31];
assign DFI_WRDATA_P2_slice_63[63]                          = DFI_WRDATA_P2[63:63];
assign DFI_WRDATA_P3_slice_0[0]                            = DFI_WRDATA_P3[0:0];
assign DFI_WRDATA_P3_slice_1[32]                           = DFI_WRDATA_P3[32:32];
assign DFI_WRDATA_P3_slice_2[1]                            = DFI_WRDATA_P3[1:1];
assign DFI_WRDATA_P3_slice_3[33]                           = DFI_WRDATA_P3[33:33];
assign DFI_WRDATA_P3_slice_4[2]                            = DFI_WRDATA_P3[2:2];
assign DFI_WRDATA_P3_slice_5[34]                           = DFI_WRDATA_P3[34:34];
assign DFI_WRDATA_P3_slice_6[3]                            = DFI_WRDATA_P3[3:3];
assign DFI_WRDATA_P3_slice_7[35]                           = DFI_WRDATA_P3[35:35];
assign DFI_WRDATA_P3_slice_8[4]                            = DFI_WRDATA_P3[4:4];
assign DFI_WRDATA_P3_slice_9[36]                           = DFI_WRDATA_P3[36:36];
assign DFI_WRDATA_P3_slice_10[5]                           = DFI_WRDATA_P3[5:5];
assign DFI_WRDATA_P3_slice_11[37]                          = DFI_WRDATA_P3[37:37];
assign DFI_WRDATA_P3_slice_12[6]                           = DFI_WRDATA_P3[6:6];
assign DFI_WRDATA_P3_slice_13[38]                          = DFI_WRDATA_P3[38:38];
assign DFI_WRDATA_P3_slice_14[7]                           = DFI_WRDATA_P3[7:7];
assign DFI_WRDATA_P3_slice_15[39]                          = DFI_WRDATA_P3[39:39];
assign DFI_WRDATA_P3_slice_16[8]                           = DFI_WRDATA_P3[8:8];
assign DFI_WRDATA_P3_slice_17[40]                          = DFI_WRDATA_P3[40:40];
assign DFI_WRDATA_P3_slice_18[9]                           = DFI_WRDATA_P3[9:9];
assign DFI_WRDATA_P3_slice_19[41]                          = DFI_WRDATA_P3[41:41];
assign DFI_WRDATA_P3_slice_20[10]                          = DFI_WRDATA_P3[10:10];
assign DFI_WRDATA_P3_slice_21[42]                          = DFI_WRDATA_P3[42:42];
assign DFI_WRDATA_P3_slice_22[11]                          = DFI_WRDATA_P3[11:11];
assign DFI_WRDATA_P3_slice_23[43]                          = DFI_WRDATA_P3[43:43];
assign DFI_WRDATA_P3_slice_24[12]                          = DFI_WRDATA_P3[12:12];
assign DFI_WRDATA_P3_slice_25[44]                          = DFI_WRDATA_P3[44:44];
assign DFI_WRDATA_P3_slice_26[13]                          = DFI_WRDATA_P3[13:13];
assign DFI_WRDATA_P3_slice_27[45]                          = DFI_WRDATA_P3[45:45];
assign DFI_WRDATA_P3_slice_28[14]                          = DFI_WRDATA_P3[14:14];
assign DFI_WRDATA_P3_slice_29[46]                          = DFI_WRDATA_P3[46:46];
assign DFI_WRDATA_P3_slice_30[15]                          = DFI_WRDATA_P3[15:15];
assign DFI_WRDATA_P3_slice_31[47]                          = DFI_WRDATA_P3[47:47];
assign DFI_WRDATA_P3_slice_32[16]                          = DFI_WRDATA_P3[16:16];
assign DFI_WRDATA_P3_slice_33[48]                          = DFI_WRDATA_P3[48:48];
assign DFI_WRDATA_P3_slice_34[17]                          = DFI_WRDATA_P3[17:17];
assign DFI_WRDATA_P3_slice_35[49]                          = DFI_WRDATA_P3[49:49];
assign DFI_WRDATA_P3_slice_36[18]                          = DFI_WRDATA_P3[18:18];
assign DFI_WRDATA_P3_slice_37[50]                          = DFI_WRDATA_P3[50:50];
assign DFI_WRDATA_P3_slice_38[19]                          = DFI_WRDATA_P3[19:19];
assign DFI_WRDATA_P3_slice_39[51]                          = DFI_WRDATA_P3[51:51];
assign DFI_WRDATA_P3_slice_40[20]                          = DFI_WRDATA_P3[20:20];
assign DFI_WRDATA_P3_slice_41[52]                          = DFI_WRDATA_P3[52:52];
assign DFI_WRDATA_P3_slice_42[21]                          = DFI_WRDATA_P3[21:21];
assign DFI_WRDATA_P3_slice_43[53]                          = DFI_WRDATA_P3[53:53];
assign DFI_WRDATA_P3_slice_44[22]                          = DFI_WRDATA_P3[22:22];
assign DFI_WRDATA_P3_slice_45[54]                          = DFI_WRDATA_P3[54:54];
assign DFI_WRDATA_P3_slice_46[23]                          = DFI_WRDATA_P3[23:23];
assign DFI_WRDATA_P3_slice_47[55]                          = DFI_WRDATA_P3[55:55];
assign DFI_WRDATA_P3_slice_48[24]                          = DFI_WRDATA_P3[24:24];
assign DFI_WRDATA_P3_slice_49[56]                          = DFI_WRDATA_P3[56:56];
assign DFI_WRDATA_P3_slice_50[25]                          = DFI_WRDATA_P3[25:25];
assign DFI_WRDATA_P3_slice_51[57]                          = DFI_WRDATA_P3[57:57];
assign DFI_WRDATA_P3_slice_52[26]                          = DFI_WRDATA_P3[26:26];
assign DFI_WRDATA_P3_slice_53[58]                          = DFI_WRDATA_P3[58:58];
assign DFI_WRDATA_P3_slice_54[27]                          = DFI_WRDATA_P3[27:27];
assign DFI_WRDATA_P3_slice_55[59]                          = DFI_WRDATA_P3[59:59];
assign DFI_WRDATA_P3_slice_56[28]                          = DFI_WRDATA_P3[28:28];
assign DFI_WRDATA_P3_slice_57[60]                          = DFI_WRDATA_P3[60:60];
assign DFI_WRDATA_P3_slice_58[29]                          = DFI_WRDATA_P3[29:29];
assign DFI_WRDATA_P3_slice_59[61]                          = DFI_WRDATA_P3[61:61];
assign DFI_WRDATA_P3_slice_60[30]                          = DFI_WRDATA_P3[30:30];
assign DFI_WRDATA_P3_slice_61[62]                          = DFI_WRDATA_P3[62:62];
assign DFI_WRDATA_P3_slice_62[31]                          = DFI_WRDATA_P3[31:31];
assign DFI_WRDATA_P3_slice_63[63]                          = DFI_WRDATA_P3[63:63];
assign IOD_A_12_RX_DATA_03to3[3]                           = RX_DATA_0_net_0[3:3];
assign IOD_BCLK_TRAINING_RX_DATA_00to0[0]                  = RX_DATA_0_net_1[0:0];
assign IOD_BCLK_TRAINING_RX_DATA_02to2[2]                  = RX_DATA_0_net_1[2:2];
assign IOD_BCLK_TRAINING_RX_DATA_04to4[4]                  = RX_DATA_0_net_1[4:4];
assign IOD_BCLK_TRAINING_RX_DATA_06to6[6]                  = RX_DATA_0_net_1[6:6];
assign IOD_REF_CLK_TRAINING_RX_DATA_06to6[6]               = RX_DATA_0_net_2[6:6];
assign IOD_TRAINING_0_CLK_SEL0to0[0]                       = CLK_SEL_net_0[0:0];
assign IOD_TRAINING_0_CLK_SEL1to1[1]                       = CLK_SEL_net_0[1:1];
assign IOD_TRAINING_0_CLK_SEL2to2[2]                       = CLK_SEL_net_0[2:2];
assign IOD_TRAINING_0_CLK_SEL3to3[3]                       = CLK_SEL_net_0[3:3];
assign IOD_TRAINING_0_CLK_SEL4to4[4]                       = CLK_SEL_net_0[4:4];
assign IOD_TRAINING_0_CLK_SEL5to5[5]                       = CLK_SEL_net_0[5:5];
assign IOD_TRAINING_0_CLK_SEL6to6[6]                       = CLK_SEL_net_0[6:6];
assign IOD_TRAINING_0_CLK_SEL7to7[7]                       = CLK_SEL_net_0[7:7];
assign IOD_TRAINING_0_CLK_SEL8to8[8]                       = CLK_SEL_net_0[8:8];
assign IOD_TRAINING_0_CLK_SEL9to9[9]                       = CLK_SEL_net_0[9:9];
assign IOD_TRAINING_0_CLK_SEL10to10[10]                    = CLK_SEL_net_0[10:10];
assign IOD_TRAINING_0_CLK_SEL11to11[11]                    = CLK_SEL_net_0[11:11];
assign IOD_TRAINING_0_DELAY_LINE_SEL_RD0to0[0]             = DELAY_LINE_SEL_RD_net_0[0:0];
assign IOD_TRAINING_0_DELAY_LINE_SEL_RD1to1[1]             = DELAY_LINE_SEL_RD_net_0[1:1];
assign IOD_TRAINING_0_DELAY_LINE_SEL_RD2to2[2]             = DELAY_LINE_SEL_RD_net_0[2:2];
assign IOD_TRAINING_0_DELAY_LINE_SEL_RD3to3[3]             = DELAY_LINE_SEL_RD_net_0[3:3];
assign IOD_TRAINING_0_DFI_BANK_P0_OUT0to0[0]               = DFI_BANK_P0_OUT_net_0[0:0];
assign IOD_TRAINING_0_DFI_BANK_P0_OUT1to1[1]               = DFI_BANK_P0_OUT_net_0[1:1];
assign IOD_TRAINING_0_DFI_BANK_P1_OUT0to0[0]               = DFI_BANK_P1_OUT_net_0[0:0];
assign IOD_TRAINING_0_DFI_BANK_P1_OUT1to1[1]               = DFI_BANK_P1_OUT_net_0[1:1];
assign IOD_TRAINING_0_DFI_BANK_P2_OUT0to0[0]               = DFI_BANK_P2_OUT_net_0[0:0];
assign IOD_TRAINING_0_DFI_BANK_P2_OUT1to1[1]               = DFI_BANK_P2_OUT_net_0[1:1];
assign IOD_TRAINING_0_DFI_BANK_P3_OUT0to0[0]               = DFI_BANK_P3_OUT_net_0[0:0];
assign IOD_TRAINING_0_DFI_BANK_P3_OUT1to1[1]               = DFI_BANK_P3_OUT_net_0[1:1];
assign IOD_TRAINING_0_DFI_BG_P0_OUT0to0[0]                 = DFI_BG_P0_OUT_net_0[0:0];
assign IOD_TRAINING_0_DFI_BG_P0_OUT1to1[1]                 = DFI_BG_P0_OUT_net_0[1:1];
assign IOD_TRAINING_0_DFI_BG_P1_OUT0to0[0]                 = DFI_BG_P1_OUT_net_0[0:0];
assign IOD_TRAINING_0_DFI_BG_P1_OUT1to1[1]                 = DFI_BG_P1_OUT_net_0[1:1];
assign IOD_TRAINING_0_DFI_BG_P2_OUT0to0[0]                 = DFI_BG_P2_OUT_net_0[0:0];
assign IOD_TRAINING_0_DFI_BG_P2_OUT1to1[1]                 = DFI_BG_P2_OUT_net_0[1:1];
assign IOD_TRAINING_0_DFI_BG_P3_OUT0to0[0]                 = DFI_BG_P3_OUT_net_0[0:0];
assign IOD_TRAINING_0_DFI_BG_P3_OUT1to1[1]                 = DFI_BG_P3_OUT_net_0[1:1];
assign IOD_TRAINING_0_DIRECTION0to0[0]                     = DIRECTION_net_0[0:0];
assign IOD_TRAINING_0_DIRECTION1to1[1]                     = DIRECTION_net_0[1:1];
assign IOD_TRAINING_0_DIRECTION2to2[2]                     = DIRECTION_net_0[2:2];
assign IOD_TRAINING_0_DIRECTION3to3[3]                     = DIRECTION_net_0[3:3];
assign IOD_TRAINING_0_DIRECTION4to4[4]                     = DIRECTION_net_0[4:4];
assign IOD_TRAINING_0_DIRECTION5to5[5]                     = DIRECTION_net_0[5:5];
assign IOD_TRAINING_0_DIRECTION6to6[6]                     = DIRECTION_net_0[6:6];
assign IOD_TRAINING_0_DIRECTION7to7[7]                     = DIRECTION_net_0[7:7];
assign IOD_TRAINING_0_DIRECTION8to8[8]                     = DIRECTION_net_0[8:8];
assign IOD_TRAINING_0_DIRECTION9to9[9]                     = DIRECTION_net_0[9:9];
assign IOD_TRAINING_0_DIRECTION10to10[10]                  = DIRECTION_net_0[10:10];
assign IOD_TRAINING_0_DIRECTION11to11[11]                  = DIRECTION_net_0[11:11];
assign IOD_TRAINING_0_DIRECTION12to12[12]                  = DIRECTION_net_0[12:12];
assign IOD_TRAINING_0_DIRECTION13to13[13]                  = DIRECTION_net_0[13:13];
assign IOD_TRAINING_0_DIRECTION14to14[14]                  = DIRECTION_net_0[14:14];
assign IOD_TRAINING_0_DIRECTION15to15[15]                  = DIRECTION_net_0[15:15];
assign IOD_TRAINING_0_DIRECTION16to16[16]                  = DIRECTION_net_0[16:16];
assign IOD_TRAINING_0_DIRECTION17to17[17]                  = DIRECTION_net_0[17:17];
assign IOD_TRAINING_0_DIRECTION18to18[18]                  = DIRECTION_net_0[18:18];
assign IOD_TRAINING_0_DIRECTION19to19[19]                  = DIRECTION_net_0[19:19];
assign IOD_TRAINING_0_DIRECTION20to20[20]                  = DIRECTION_net_0[20:20];
assign IOD_TRAINING_0_DIRECTION21to21[21]                  = DIRECTION_net_0[21:21];
assign IOD_TRAINING_0_DIRECTION22to22[22]                  = DIRECTION_net_0[22:22];
assign IOD_TRAINING_0_DIRECTION23to23[23]                  = DIRECTION_net_0[23:23];
assign IOD_TRAINING_0_DIRECTION24to24[24]                  = DIRECTION_net_0[24:24];
assign IOD_TRAINING_0_DIRECTION25to25[25]                  = DIRECTION_net_0[25:25];
assign IOD_TRAINING_0_DIRECTION26to26[26]                  = DIRECTION_net_0[26:26];
assign IOD_TRAINING_0_DIRECTION27to27[27]                  = DIRECTION_net_0[27:27];
assign IOD_TRAINING_0_DIRECTION28to28[28]                  = DIRECTION_net_0[28:28];
assign IOD_TRAINING_0_DIRECTION29to29[29]                  = DIRECTION_net_0[29:29];
assign IOD_TRAINING_0_DIRECTION30to30[30]                  = DIRECTION_net_0[30:30];
assign IOD_TRAINING_0_DIRECTION31to31[31]                  = DIRECTION_net_0[31:31];
assign IOD_TRAINING_0_DIRECTION32to32[32]                  = DIRECTION_net_0[32:32];
assign IOD_TRAINING_0_DIRECTION33to33[33]                  = DIRECTION_net_0[33:33];
assign IOD_TRAINING_0_DIRECTION34to34[34]                  = DIRECTION_net_0[34:34];
assign IOD_TRAINING_0_DIRECTION35to35[35]                  = DIRECTION_net_0[35:35];
assign IOD_TRAINING_0_DM_OE_P00to0[0]                      = DM_OE_P0_net_0[0:0];
assign IOD_TRAINING_0_DM_OE_P01to1[1]                      = DM_OE_P0_net_0[1:1];
assign IOD_TRAINING_0_DM_OE_P02to2[2]                      = DM_OE_P0_net_0[2:2];
assign IOD_TRAINING_0_DM_OE_P03to3[3]                      = DM_OE_P0_net_0[3:3];
assign IOD_TRAINING_0_DM_OE_P10to0[0]                      = DM_OE_P1_net_0[0:0];
assign IOD_TRAINING_0_DM_OE_P11to1[1]                      = DM_OE_P1_net_0[1:1];
assign IOD_TRAINING_0_DM_OE_P12to2[2]                      = DM_OE_P1_net_0[2:2];
assign IOD_TRAINING_0_DM_OE_P13to3[3]                      = DM_OE_P1_net_0[3:3];
assign IOD_TRAINING_0_DM_OE_P20to0[0]                      = DM_OE_P2_net_0[0:0];
assign IOD_TRAINING_0_DM_OE_P21to1[1]                      = DM_OE_P2_net_0[1:1];
assign IOD_TRAINING_0_DM_OE_P22to2[2]                      = DM_OE_P2_net_0[2:2];
assign IOD_TRAINING_0_DM_OE_P23to3[3]                      = DM_OE_P2_net_0[3:3];
assign IOD_TRAINING_0_DM_OE_P30to0[0]                      = DM_OE_P3_net_0[0:0];
assign IOD_TRAINING_0_DM_OE_P31to1[1]                      = DM_OE_P3_net_0[1:1];
assign IOD_TRAINING_0_DM_OE_P32to2[2]                      = DM_OE_P3_net_0[2:2];
assign IOD_TRAINING_0_DM_OE_P33to3[3]                      = DM_OE_P3_net_0[3:3];
assign IOD_TRAINING_0_DQS_OE_P00to0[0]                     = DQS_OE_P0_net_0[0:0];
assign IOD_TRAINING_0_DQS_OE_P01to1[1]                     = DQS_OE_P0_net_0[1:1];
assign IOD_TRAINING_0_DQS_OE_P02to2[2]                     = DQS_OE_P0_net_0[2:2];
assign IOD_TRAINING_0_DQS_OE_P03to3[3]                     = DQS_OE_P0_net_0[3:3];
assign IOD_TRAINING_0_DQS_OE_P10to0[0]                     = DQS_OE_P1_net_0[0:0];
assign IOD_TRAINING_0_DQS_OE_P11to1[1]                     = DQS_OE_P1_net_0[1:1];
assign IOD_TRAINING_0_DQS_OE_P12to2[2]                     = DQS_OE_P1_net_0[2:2];
assign IOD_TRAINING_0_DQS_OE_P13to3[3]                     = DQS_OE_P1_net_0[3:3];
assign IOD_TRAINING_0_DQS_OE_P20to0[0]                     = DQS_OE_P2_net_0[0:0];
assign IOD_TRAINING_0_DQS_OE_P21to1[1]                     = DQS_OE_P2_net_0[1:1];
assign IOD_TRAINING_0_DQS_OE_P22to2[2]                     = DQS_OE_P2_net_0[2:2];
assign IOD_TRAINING_0_DQS_OE_P23to3[3]                     = DQS_OE_P2_net_0[3:3];
assign IOD_TRAINING_0_DQS_OE_P30to0[0]                     = DQS_OE_P3_net_0[0:0];
assign IOD_TRAINING_0_DQS_OE_P31to1[1]                     = DQS_OE_P3_net_0[1:1];
assign IOD_TRAINING_0_DQS_OE_P32to2[2]                     = DQS_OE_P3_net_0[2:2];
assign IOD_TRAINING_0_DQS_OE_P33to3[3]                     = DQS_OE_P3_net_0[3:3];
assign IOD_TRAINING_0_DQSW270_DELAY_LINE_DIRECTION0to0[0]  = DQSW270_DELAY_LINE_DIRECTION_net_0[0:0];
assign IOD_TRAINING_0_DQSW270_DELAY_LINE_DIRECTION1to1[1]  = DQSW270_DELAY_LINE_DIRECTION_net_0[1:1];
assign IOD_TRAINING_0_DQSW270_DELAY_LINE_DIRECTION2to2[2]  = DQSW270_DELAY_LINE_DIRECTION_net_0[2:2];
assign IOD_TRAINING_0_DQSW270_DELAY_LINE_DIRECTION3to3[3]  = DQSW270_DELAY_LINE_DIRECTION_net_0[3:3];
assign IOD_TRAINING_0_DQSW270_DELAY_LINE_LOAD0to0[0]       = DQSW270_DELAY_LINE_LOAD_net_0[0:0];
assign IOD_TRAINING_0_DQSW270_DELAY_LINE_LOAD1to1[1]       = DQSW270_DELAY_LINE_LOAD_net_0[1:1];
assign IOD_TRAINING_0_DQSW270_DELAY_LINE_LOAD2to2[2]       = DQSW270_DELAY_LINE_LOAD_net_0[2:2];
assign IOD_TRAINING_0_DQSW270_DELAY_LINE_LOAD3to3[3]       = DQSW270_DELAY_LINE_LOAD_net_0[3:3];
assign IOD_TRAINING_0_DQSW270_DELAY_LINE_MOVE0to0[0]       = DQSW270_DELAY_LINE_MOVE_net_0[0:0];
assign IOD_TRAINING_0_DQSW270_DELAY_LINE_MOVE1to1[1]       = DQSW270_DELAY_LINE_MOVE_net_0[1:1];
assign IOD_TRAINING_0_DQSW270_DELAY_LINE_MOVE2to2[2]       = DQSW270_DELAY_LINE_MOVE_net_0[2:2];
assign IOD_TRAINING_0_DQSW270_DELAY_LINE_MOVE3to3[3]       = DQSW270_DELAY_LINE_MOVE_net_0[3:3];
assign IOD_TRAINING_0_DQSW270_EYE_MONITOR_CLR_FLAGS0to0[0] = DQSW270_EYE_MONITOR_CLR_FLAGS_net_0[0:0];
assign IOD_TRAINING_0_DQSW270_EYE_MONITOR_CLR_FLAGS1to1[1] = DQSW270_EYE_MONITOR_CLR_FLAGS_net_0[1:1];
assign IOD_TRAINING_0_DQSW270_EYE_MONITOR_CLR_FLAGS2to2[2] = DQSW270_EYE_MONITOR_CLR_FLAGS_net_0[2:2];
assign IOD_TRAINING_0_DQSW270_EYE_MONITOR_CLR_FLAGS3to3[3] = DQSW270_EYE_MONITOR_CLR_FLAGS_net_0[3:3];
assign IOD_TRAINING_0_DQSW_DELAY_LINE_DIRECTION0to0[0]     = DQSW_DELAY_LINE_DIRECTION_net_0[0:0];
assign IOD_TRAINING_0_DQSW_DELAY_LINE_DIRECTION1to1[1]     = DQSW_DELAY_LINE_DIRECTION_net_0[1:1];
assign IOD_TRAINING_0_DQSW_DELAY_LINE_DIRECTION2to2[2]     = DQSW_DELAY_LINE_DIRECTION_net_0[2:2];
assign IOD_TRAINING_0_DQSW_DELAY_LINE_DIRECTION3to3[3]     = DQSW_DELAY_LINE_DIRECTION_net_0[3:3];
assign IOD_TRAINING_0_DQSW_DELAY_LINE_LOAD0to0[0]          = DQSW_DELAY_LINE_LOAD_net_0[0:0];
assign IOD_TRAINING_0_DQSW_DELAY_LINE_LOAD1to1[1]          = DQSW_DELAY_LINE_LOAD_net_0[1:1];
assign IOD_TRAINING_0_DQSW_DELAY_LINE_LOAD2to2[2]          = DQSW_DELAY_LINE_LOAD_net_0[2:2];
assign IOD_TRAINING_0_DQSW_DELAY_LINE_LOAD3to3[3]          = DQSW_DELAY_LINE_LOAD_net_0[3:3];
assign IOD_TRAINING_0_DQSW_DELAY_LINE_MOVE0to0[0]          = DQSW_DELAY_LINE_MOVE_net_0[0:0];
assign IOD_TRAINING_0_DQSW_DELAY_LINE_MOVE1to1[1]          = DQSW_DELAY_LINE_MOVE_net_0[1:1];
assign IOD_TRAINING_0_DQSW_DELAY_LINE_MOVE2to2[2]          = DQSW_DELAY_LINE_MOVE_net_0[2:2];
assign IOD_TRAINING_0_DQSW_DELAY_LINE_MOVE3to3[3]          = DQSW_DELAY_LINE_MOVE_net_0[3:3];
assign IOD_TRAINING_0_DQSW_EYE_MONITOR_CLR_FLAGS0to0[0]    = DQSW_EYE_MONITOR_CLR_FLAGS_net_0[0:0];
assign IOD_TRAINING_0_DQSW_EYE_MONITOR_CLR_FLAGS1to1[1]    = DQSW_EYE_MONITOR_CLR_FLAGS_net_0[1:1];
assign IOD_TRAINING_0_DQSW_EYE_MONITOR_CLR_FLAGS2to2[2]    = DQSW_EYE_MONITOR_CLR_FLAGS_net_0[2:2];
assign IOD_TRAINING_0_DQSW_EYE_MONITOR_CLR_FLAGS3to3[3]    = DQSW_EYE_MONITOR_CLR_FLAGS_net_0[3:3];
assign IOD_TRAINING_0_DQSW_SELA7to0                        = DQSW_SELA_net_0[7:0];
assign IOD_TRAINING_0_DQSW_SELA15to8                       = DQSW_SELA_net_0[15:8];
assign IOD_TRAINING_0_DQSW_SELA23to16                      = DQSW_SELA_net_0[23:16];
assign IOD_TRAINING_0_DQSW_SELA31to24                      = DQSW_SELA_net_0[31:24];
assign IOD_TRAINING_0_INIT_PAUSE0to0[0]                    = INIT_PAUSE_net_0[0:0];
assign IOD_TRAINING_0_INIT_PAUSE1to1[1]                    = INIT_PAUSE_net_0[1:1];
assign IOD_TRAINING_0_INIT_PAUSE2to2[2]                    = INIT_PAUSE_net_0[2:2];
assign IOD_TRAINING_0_INIT_PAUSE3to3[3]                    = INIT_PAUSE_net_0[3:3];
assign IOD_TRAINING_0_IOG_ADDRESS_P00to0[0]                = IOG_ADDRESS_P0_net_0[0:0];
assign IOD_TRAINING_0_IOG_ADDRESS_P01to1[1]                = IOG_ADDRESS_P0_net_0[1:1];
assign IOD_TRAINING_0_IOG_ADDRESS_P02to2[2]                = IOG_ADDRESS_P0_net_0[2:2];
assign IOD_TRAINING_0_IOG_ADDRESS_P03to3[3]                = IOG_ADDRESS_P0_net_0[3:3];
assign IOD_TRAINING_0_IOG_ADDRESS_P04to4[4]                = IOG_ADDRESS_P0_net_0[4:4];
assign IOD_TRAINING_0_IOG_ADDRESS_P05to5[5]                = IOG_ADDRESS_P0_net_0[5:5];
assign IOD_TRAINING_0_IOG_ADDRESS_P06to6[6]                = IOG_ADDRESS_P0_net_0[6:6];
assign IOD_TRAINING_0_IOG_ADDRESS_P07to7[7]                = IOG_ADDRESS_P0_net_0[7:7];
assign IOD_TRAINING_0_IOG_ADDRESS_P08to8[8]                = IOG_ADDRESS_P0_net_0[8:8];
assign IOD_TRAINING_0_IOG_ADDRESS_P09to9[9]                = IOG_ADDRESS_P0_net_0[9:9];
assign IOD_TRAINING_0_IOG_ADDRESS_P10to0[0]                = IOG_ADDRESS_P1_net_0[0:0];
assign IOD_TRAINING_0_IOG_ADDRESS_P010to10[10]             = IOG_ADDRESS_P0_net_0[10:10];
assign IOD_TRAINING_0_IOG_ADDRESS_P11to1[1]                = IOG_ADDRESS_P1_net_0[1:1];
assign IOD_TRAINING_0_IOG_ADDRESS_P011to11[11]             = IOG_ADDRESS_P0_net_0[11:11];
assign IOD_TRAINING_0_IOG_ADDRESS_P12to2[2]                = IOG_ADDRESS_P1_net_0[2:2];
assign IOD_TRAINING_0_IOG_ADDRESS_P012to12[12]             = IOG_ADDRESS_P0_net_0[12:12];
assign IOD_TRAINING_0_IOG_ADDRESS_P13to3[3]                = IOG_ADDRESS_P1_net_0[3:3];
assign IOD_TRAINING_0_IOG_ADDRESS_P013to13[13]             = IOG_ADDRESS_P0_net_0[13:13];
assign IOD_TRAINING_0_IOG_ADDRESS_P14to4[4]                = IOG_ADDRESS_P1_net_0[4:4];
assign IOD_TRAINING_0_IOG_ADDRESS_P15to5[5]                = IOG_ADDRESS_P1_net_0[5:5];
assign IOD_TRAINING_0_IOG_ADDRESS_P16to6[6]                = IOG_ADDRESS_P1_net_0[6:6];
assign IOD_TRAINING_0_IOG_ADDRESS_P17to7[7]                = IOG_ADDRESS_P1_net_0[7:7];
assign IOD_TRAINING_0_IOG_ADDRESS_P18to8[8]                = IOG_ADDRESS_P1_net_0[8:8];
assign IOD_TRAINING_0_IOG_ADDRESS_P19to9[9]                = IOG_ADDRESS_P1_net_0[9:9];
assign IOD_TRAINING_0_IOG_ADDRESS_P20to0[0]                = IOG_ADDRESS_P2_net_0[0:0];
assign IOD_TRAINING_0_IOG_ADDRESS_P21to1[1]                = IOG_ADDRESS_P2_net_0[1:1];
assign IOD_TRAINING_0_IOG_ADDRESS_P22to2[2]                = IOG_ADDRESS_P2_net_0[2:2];
assign IOD_TRAINING_0_IOG_ADDRESS_P23to3[3]                = IOG_ADDRESS_P2_net_0[3:3];
assign IOD_TRAINING_0_IOG_ADDRESS_P24to4[4]                = IOG_ADDRESS_P2_net_0[4:4];
assign IOD_TRAINING_0_IOG_ADDRESS_P25to5[5]                = IOG_ADDRESS_P2_net_0[5:5];
assign IOD_TRAINING_0_IOG_ADDRESS_P26to6[6]                = IOG_ADDRESS_P2_net_0[6:6];
assign IOD_TRAINING_0_IOG_ADDRESS_P27to7[7]                = IOG_ADDRESS_P2_net_0[7:7];
assign IOD_TRAINING_0_IOG_ADDRESS_P28to8[8]                = IOG_ADDRESS_P2_net_0[8:8];
assign IOD_TRAINING_0_IOG_ADDRESS_P29to9[9]                = IOG_ADDRESS_P2_net_0[9:9];
assign IOD_TRAINING_0_IOG_ADDRESS_P30to0[0]                = IOG_ADDRESS_P3_net_0[0:0];
assign IOD_TRAINING_0_IOG_ADDRESS_P31to1[1]                = IOG_ADDRESS_P3_net_0[1:1];
assign IOD_TRAINING_0_IOG_ADDRESS_P32to2[2]                = IOG_ADDRESS_P3_net_0[2:2];
assign IOD_TRAINING_0_IOG_ADDRESS_P33to3[3]                = IOG_ADDRESS_P3_net_0[3:3];
assign IOD_TRAINING_0_IOG_ADDRESS_P34to4[4]                = IOG_ADDRESS_P3_net_0[4:4];
assign IOD_TRAINING_0_IOG_ADDRESS_P35to5[5]                = IOG_ADDRESS_P3_net_0[5:5];
assign IOD_TRAINING_0_IOG_ADDRESS_P36to6[6]                = IOG_ADDRESS_P3_net_0[6:6];
assign IOD_TRAINING_0_IOG_ADDRESS_P37to7[7]                = IOG_ADDRESS_P3_net_0[7:7];
assign IOD_TRAINING_0_IOG_ADDRESS_P38to8[8]                = IOG_ADDRESS_P3_net_0[8:8];
assign IOD_TRAINING_0_IOG_ADDRESS_P39to9[9]                = IOG_ADDRESS_P3_net_0[9:9];
assign IOD_TRAINING_0_IOG_ADDRESS_P110to10[10]             = IOG_ADDRESS_P1_net_0[10:10];
assign IOD_TRAINING_0_IOG_ADDRESS_P111to11[11]             = IOG_ADDRESS_P1_net_0[11:11];
assign IOD_TRAINING_0_IOG_ADDRESS_P112to12[12]             = IOG_ADDRESS_P1_net_0[12:12];
assign IOD_TRAINING_0_IOG_ADDRESS_P113to13[13]             = IOG_ADDRESS_P1_net_0[13:13];
assign IOD_TRAINING_0_IOG_ADDRESS_P210to10[10]             = IOG_ADDRESS_P2_net_0[10:10];
assign IOD_TRAINING_0_IOG_ADDRESS_P211to11[11]             = IOG_ADDRESS_P2_net_0[11:11];
assign IOD_TRAINING_0_IOG_ADDRESS_P212to12[12]             = IOG_ADDRESS_P2_net_0[12:12];
assign IOD_TRAINING_0_IOG_ADDRESS_P213to13[13]             = IOG_ADDRESS_P2_net_0[13:13];
assign IOD_TRAINING_0_IOG_ADDRESS_P310to10[10]             = IOG_ADDRESS_P3_net_0[10:10];
assign IOD_TRAINING_0_IOG_ADDRESS_P311to11[11]             = IOG_ADDRESS_P3_net_0[11:11];
assign IOD_TRAINING_0_IOG_ADDRESS_P312to12[12]             = IOG_ADDRESS_P3_net_0[12:12];
assign IOD_TRAINING_0_IOG_ADDRESS_P313to13[13]             = IOG_ADDRESS_P3_net_0[13:13];
assign IOD_TRAINING_0_IOG_DM_TXDATA_OUT0to0[0]             = IOG_DM_TXDATA_OUT_net_0[0:0];
assign IOD_TRAINING_0_IOG_DM_TXDATA_OUT1to1[1]             = IOG_DM_TXDATA_OUT_net_0[1:1];
assign IOD_TRAINING_0_IOG_DM_TXDATA_OUT2to2[2]             = IOG_DM_TXDATA_OUT_net_0[2:2];
assign IOD_TRAINING_0_IOG_DM_TXDATA_OUT3to3[3]             = IOG_DM_TXDATA_OUT_net_0[3:3];
assign IOD_TRAINING_0_IOG_DM_TXDATA_OUT4to4[4]             = IOG_DM_TXDATA_OUT_net_0[4:4];
assign IOD_TRAINING_0_IOG_DM_TXDATA_OUT5to5[5]             = IOG_DM_TXDATA_OUT_net_0[5:5];
assign IOD_TRAINING_0_IOG_DM_TXDATA_OUT6to6[6]             = IOG_DM_TXDATA_OUT_net_0[6:6];
assign IOD_TRAINING_0_IOG_DM_TXDATA_OUT7to7[7]             = IOG_DM_TXDATA_OUT_net_0[7:7];
assign IOD_TRAINING_0_IOG_DM_TXDATA_OUT8to8[8]             = IOG_DM_TXDATA_OUT_net_0[8:8];
assign IOD_TRAINING_0_IOG_DM_TXDATA_OUT9to9[9]             = IOG_DM_TXDATA_OUT_net_0[9:9];
assign IOD_TRAINING_0_IOG_DM_TXDATA_OUT10to10[10]          = IOG_DM_TXDATA_OUT_net_0[10:10];
assign IOD_TRAINING_0_IOG_DM_TXDATA_OUT11to11[11]          = IOG_DM_TXDATA_OUT_net_0[11:11];
assign IOD_TRAINING_0_IOG_DM_TXDATA_OUT12to12[12]          = IOG_DM_TXDATA_OUT_net_0[12:12];
assign IOD_TRAINING_0_IOG_DM_TXDATA_OUT13to13[13]          = IOG_DM_TXDATA_OUT_net_0[13:13];
assign IOD_TRAINING_0_IOG_DM_TXDATA_OUT14to14[14]          = IOG_DM_TXDATA_OUT_net_0[14:14];
assign IOD_TRAINING_0_IOG_DM_TXDATA_OUT15to15[15]          = IOG_DM_TXDATA_OUT_net_0[15:15];
assign IOD_TRAINING_0_IOG_DM_TXDATA_OUT16to16[16]          = IOG_DM_TXDATA_OUT_net_0[16:16];
assign IOD_TRAINING_0_IOG_DM_TXDATA_OUT17to17[17]          = IOG_DM_TXDATA_OUT_net_0[17:17];
assign IOD_TRAINING_0_IOG_DM_TXDATA_OUT18to18[18]          = IOG_DM_TXDATA_OUT_net_0[18:18];
assign IOD_TRAINING_0_IOG_DM_TXDATA_OUT19to19[19]          = IOG_DM_TXDATA_OUT_net_0[19:19];
assign IOD_TRAINING_0_IOG_DM_TXDATA_OUT20to20[20]          = IOG_DM_TXDATA_OUT_net_0[20:20];
assign IOD_TRAINING_0_IOG_DM_TXDATA_OUT21to21[21]          = IOG_DM_TXDATA_OUT_net_0[21:21];
assign IOD_TRAINING_0_IOG_DM_TXDATA_OUT22to22[22]          = IOG_DM_TXDATA_OUT_net_0[22:22];
assign IOD_TRAINING_0_IOG_DM_TXDATA_OUT23to23[23]          = IOG_DM_TXDATA_OUT_net_0[23:23];
assign IOD_TRAINING_0_IOG_DM_TXDATA_OUT24to24[24]          = IOG_DM_TXDATA_OUT_net_0[24:24];
assign IOD_TRAINING_0_IOG_DM_TXDATA_OUT25to25[25]          = IOG_DM_TXDATA_OUT_net_0[25:25];
assign IOD_TRAINING_0_IOG_DM_TXDATA_OUT26to26[26]          = IOG_DM_TXDATA_OUT_net_0[26:26];
assign IOD_TRAINING_0_IOG_DM_TXDATA_OUT27to27[27]          = IOG_DM_TXDATA_OUT_net_0[27:27];
assign IOD_TRAINING_0_IOG_DM_TXDATA_OUT28to28[28]          = IOG_DM_TXDATA_OUT_net_0[28:28];
assign IOD_TRAINING_0_IOG_DM_TXDATA_OUT29to29[29]          = IOG_DM_TXDATA_OUT_net_0[29:29];
assign IOD_TRAINING_0_IOG_DM_TXDATA_OUT30to30[30]          = IOG_DM_TXDATA_OUT_net_0[30:30];
assign IOD_TRAINING_0_IOG_DM_TXDATA_OUT31to31[31]          = IOG_DM_TXDATA_OUT_net_0[31:31];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT0to0[0]             = IOG_DQ_TXDATA_OUT_net_0[0:0];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT1to1[1]             = IOG_DQ_TXDATA_OUT_net_0[1:1];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT2to2[2]             = IOG_DQ_TXDATA_OUT_net_0[2:2];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT3to3[3]             = IOG_DQ_TXDATA_OUT_net_0[3:3];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT4to4[4]             = IOG_DQ_TXDATA_OUT_net_0[4:4];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT5to5[5]             = IOG_DQ_TXDATA_OUT_net_0[5:5];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT6to6[6]             = IOG_DQ_TXDATA_OUT_net_0[6:6];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT7to7[7]             = IOG_DQ_TXDATA_OUT_net_0[7:7];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT8to8[8]             = IOG_DQ_TXDATA_OUT_net_0[8:8];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT9to9[9]             = IOG_DQ_TXDATA_OUT_net_0[9:9];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT10to10[10]          = IOG_DQ_TXDATA_OUT_net_0[10:10];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT11to11[11]          = IOG_DQ_TXDATA_OUT_net_0[11:11];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT12to12[12]          = IOG_DQ_TXDATA_OUT_net_0[12:12];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT13to13[13]          = IOG_DQ_TXDATA_OUT_net_0[13:13];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT14to14[14]          = IOG_DQ_TXDATA_OUT_net_0[14:14];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT15to15[15]          = IOG_DQ_TXDATA_OUT_net_0[15:15];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT16to16[16]          = IOG_DQ_TXDATA_OUT_net_0[16:16];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT17to17[17]          = IOG_DQ_TXDATA_OUT_net_0[17:17];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT18to18[18]          = IOG_DQ_TXDATA_OUT_net_0[18:18];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT19to19[19]          = IOG_DQ_TXDATA_OUT_net_0[19:19];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT20to20[20]          = IOG_DQ_TXDATA_OUT_net_0[20:20];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT21to21[21]          = IOG_DQ_TXDATA_OUT_net_0[21:21];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT22to22[22]          = IOG_DQ_TXDATA_OUT_net_0[22:22];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT23to23[23]          = IOG_DQ_TXDATA_OUT_net_0[23:23];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT24to24[24]          = IOG_DQ_TXDATA_OUT_net_0[24:24];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT25to25[25]          = IOG_DQ_TXDATA_OUT_net_0[25:25];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT26to26[26]          = IOG_DQ_TXDATA_OUT_net_0[26:26];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT27to27[27]          = IOG_DQ_TXDATA_OUT_net_0[27:27];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT28to28[28]          = IOG_DQ_TXDATA_OUT_net_0[28:28];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT29to29[29]          = IOG_DQ_TXDATA_OUT_net_0[29:29];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT30to30[30]          = IOG_DQ_TXDATA_OUT_net_0[30:30];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT31to31[31]          = IOG_DQ_TXDATA_OUT_net_0[31:31];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT32to32[32]          = IOG_DQ_TXDATA_OUT_net_0[32:32];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT33to33[33]          = IOG_DQ_TXDATA_OUT_net_0[33:33];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT34to34[34]          = IOG_DQ_TXDATA_OUT_net_0[34:34];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT35to35[35]          = IOG_DQ_TXDATA_OUT_net_0[35:35];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT36to36[36]          = IOG_DQ_TXDATA_OUT_net_0[36:36];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT37to37[37]          = IOG_DQ_TXDATA_OUT_net_0[37:37];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT38to38[38]          = IOG_DQ_TXDATA_OUT_net_0[38:38];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT39to39[39]          = IOG_DQ_TXDATA_OUT_net_0[39:39];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT40to40[40]          = IOG_DQ_TXDATA_OUT_net_0[40:40];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT41to41[41]          = IOG_DQ_TXDATA_OUT_net_0[41:41];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT42to42[42]          = IOG_DQ_TXDATA_OUT_net_0[42:42];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT43to43[43]          = IOG_DQ_TXDATA_OUT_net_0[43:43];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT44to44[44]          = IOG_DQ_TXDATA_OUT_net_0[44:44];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT45to45[45]          = IOG_DQ_TXDATA_OUT_net_0[45:45];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT46to46[46]          = IOG_DQ_TXDATA_OUT_net_0[46:46];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT47to47[47]          = IOG_DQ_TXDATA_OUT_net_0[47:47];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT48to48[48]          = IOG_DQ_TXDATA_OUT_net_0[48:48];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT49to49[49]          = IOG_DQ_TXDATA_OUT_net_0[49:49];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT50to50[50]          = IOG_DQ_TXDATA_OUT_net_0[50:50];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT51to51[51]          = IOG_DQ_TXDATA_OUT_net_0[51:51];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT52to52[52]          = IOG_DQ_TXDATA_OUT_net_0[52:52];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT53to53[53]          = IOG_DQ_TXDATA_OUT_net_0[53:53];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT54to54[54]          = IOG_DQ_TXDATA_OUT_net_0[54:54];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT55to55[55]          = IOG_DQ_TXDATA_OUT_net_0[55:55];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT56to56[56]          = IOG_DQ_TXDATA_OUT_net_0[56:56];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT57to57[57]          = IOG_DQ_TXDATA_OUT_net_0[57:57];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT58to58[58]          = IOG_DQ_TXDATA_OUT_net_0[58:58];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT59to59[59]          = IOG_DQ_TXDATA_OUT_net_0[59:59];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT60to60[60]          = IOG_DQ_TXDATA_OUT_net_0[60:60];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT61to61[61]          = IOG_DQ_TXDATA_OUT_net_0[61:61];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT62to62[62]          = IOG_DQ_TXDATA_OUT_net_0[62:62];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT63to63[63]          = IOG_DQ_TXDATA_OUT_net_0[63:63];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT64to64[64]          = IOG_DQ_TXDATA_OUT_net_0[64:64];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT65to65[65]          = IOG_DQ_TXDATA_OUT_net_0[65:65];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT66to66[66]          = IOG_DQ_TXDATA_OUT_net_0[66:66];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT67to67[67]          = IOG_DQ_TXDATA_OUT_net_0[67:67];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT68to68[68]          = IOG_DQ_TXDATA_OUT_net_0[68:68];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT69to69[69]          = IOG_DQ_TXDATA_OUT_net_0[69:69];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT70to70[70]          = IOG_DQ_TXDATA_OUT_net_0[70:70];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT71to71[71]          = IOG_DQ_TXDATA_OUT_net_0[71:71];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT72to72[72]          = IOG_DQ_TXDATA_OUT_net_0[72:72];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT73to73[73]          = IOG_DQ_TXDATA_OUT_net_0[73:73];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT74to74[74]          = IOG_DQ_TXDATA_OUT_net_0[74:74];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT75to75[75]          = IOG_DQ_TXDATA_OUT_net_0[75:75];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT76to76[76]          = IOG_DQ_TXDATA_OUT_net_0[76:76];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT77to77[77]          = IOG_DQ_TXDATA_OUT_net_0[77:77];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT78to78[78]          = IOG_DQ_TXDATA_OUT_net_0[78:78];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT79to79[79]          = IOG_DQ_TXDATA_OUT_net_0[79:79];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT80to80[80]          = IOG_DQ_TXDATA_OUT_net_0[80:80];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT81to81[81]          = IOG_DQ_TXDATA_OUT_net_0[81:81];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT82to82[82]          = IOG_DQ_TXDATA_OUT_net_0[82:82];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT83to83[83]          = IOG_DQ_TXDATA_OUT_net_0[83:83];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT84to84[84]          = IOG_DQ_TXDATA_OUT_net_0[84:84];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT85to85[85]          = IOG_DQ_TXDATA_OUT_net_0[85:85];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT86to86[86]          = IOG_DQ_TXDATA_OUT_net_0[86:86];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT87to87[87]          = IOG_DQ_TXDATA_OUT_net_0[87:87];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT88to88[88]          = IOG_DQ_TXDATA_OUT_net_0[88:88];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT89to89[89]          = IOG_DQ_TXDATA_OUT_net_0[89:89];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT90to90[90]          = IOG_DQ_TXDATA_OUT_net_0[90:90];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT91to91[91]          = IOG_DQ_TXDATA_OUT_net_0[91:91];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT92to92[92]          = IOG_DQ_TXDATA_OUT_net_0[92:92];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT93to93[93]          = IOG_DQ_TXDATA_OUT_net_0[93:93];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT94to94[94]          = IOG_DQ_TXDATA_OUT_net_0[94:94];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT95to95[95]          = IOG_DQ_TXDATA_OUT_net_0[95:95];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT96to96[96]          = IOG_DQ_TXDATA_OUT_net_0[96:96];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT97to97[97]          = IOG_DQ_TXDATA_OUT_net_0[97:97];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT98to98[98]          = IOG_DQ_TXDATA_OUT_net_0[98:98];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT99to99[99]          = IOG_DQ_TXDATA_OUT_net_0[99:99];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT100to100[100]       = IOG_DQ_TXDATA_OUT_net_0[100:100];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT101to101[101]       = IOG_DQ_TXDATA_OUT_net_0[101:101];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT102to102[102]       = IOG_DQ_TXDATA_OUT_net_0[102:102];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT103to103[103]       = IOG_DQ_TXDATA_OUT_net_0[103:103];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT104to104[104]       = IOG_DQ_TXDATA_OUT_net_0[104:104];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT105to105[105]       = IOG_DQ_TXDATA_OUT_net_0[105:105];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT106to106[106]       = IOG_DQ_TXDATA_OUT_net_0[106:106];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT107to107[107]       = IOG_DQ_TXDATA_OUT_net_0[107:107];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT108to108[108]       = IOG_DQ_TXDATA_OUT_net_0[108:108];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT109to109[109]       = IOG_DQ_TXDATA_OUT_net_0[109:109];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT110to110[110]       = IOG_DQ_TXDATA_OUT_net_0[110:110];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT111to111[111]       = IOG_DQ_TXDATA_OUT_net_0[111:111];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT112to112[112]       = IOG_DQ_TXDATA_OUT_net_0[112:112];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT113to113[113]       = IOG_DQ_TXDATA_OUT_net_0[113:113];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT114to114[114]       = IOG_DQ_TXDATA_OUT_net_0[114:114];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT115to115[115]       = IOG_DQ_TXDATA_OUT_net_0[115:115];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT116to116[116]       = IOG_DQ_TXDATA_OUT_net_0[116:116];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT117to117[117]       = IOG_DQ_TXDATA_OUT_net_0[117:117];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT118to118[118]       = IOG_DQ_TXDATA_OUT_net_0[118:118];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT119to119[119]       = IOG_DQ_TXDATA_OUT_net_0[119:119];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT120to120[120]       = IOG_DQ_TXDATA_OUT_net_0[120:120];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT121to121[121]       = IOG_DQ_TXDATA_OUT_net_0[121:121];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT122to122[122]       = IOG_DQ_TXDATA_OUT_net_0[122:122];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT123to123[123]       = IOG_DQ_TXDATA_OUT_net_0[123:123];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT124to124[124]       = IOG_DQ_TXDATA_OUT_net_0[124:124];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT125to125[125]       = IOG_DQ_TXDATA_OUT_net_0[125:125];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT126to126[126]       = IOG_DQ_TXDATA_OUT_net_0[126:126];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT127to127[127]       = IOG_DQ_TXDATA_OUT_net_0[127:127];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT128to128[128]       = IOG_DQ_TXDATA_OUT_net_0[128:128];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT129to129[129]       = IOG_DQ_TXDATA_OUT_net_0[129:129];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT130to130[130]       = IOG_DQ_TXDATA_OUT_net_0[130:130];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT131to131[131]       = IOG_DQ_TXDATA_OUT_net_0[131:131];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT132to132[132]       = IOG_DQ_TXDATA_OUT_net_0[132:132];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT133to133[133]       = IOG_DQ_TXDATA_OUT_net_0[133:133];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT134to134[134]       = IOG_DQ_TXDATA_OUT_net_0[134:134];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT135to135[135]       = IOG_DQ_TXDATA_OUT_net_0[135:135];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT136to136[136]       = IOG_DQ_TXDATA_OUT_net_0[136:136];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT137to137[137]       = IOG_DQ_TXDATA_OUT_net_0[137:137];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT138to138[138]       = IOG_DQ_TXDATA_OUT_net_0[138:138];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT139to139[139]       = IOG_DQ_TXDATA_OUT_net_0[139:139];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT140to140[140]       = IOG_DQ_TXDATA_OUT_net_0[140:140];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT141to141[141]       = IOG_DQ_TXDATA_OUT_net_0[141:141];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT142to142[142]       = IOG_DQ_TXDATA_OUT_net_0[142:142];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT143to143[143]       = IOG_DQ_TXDATA_OUT_net_0[143:143];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT144to144[144]       = IOG_DQ_TXDATA_OUT_net_0[144:144];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT145to145[145]       = IOG_DQ_TXDATA_OUT_net_0[145:145];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT146to146[146]       = IOG_DQ_TXDATA_OUT_net_0[146:146];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT147to147[147]       = IOG_DQ_TXDATA_OUT_net_0[147:147];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT148to148[148]       = IOG_DQ_TXDATA_OUT_net_0[148:148];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT149to149[149]       = IOG_DQ_TXDATA_OUT_net_0[149:149];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT150to150[150]       = IOG_DQ_TXDATA_OUT_net_0[150:150];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT151to151[151]       = IOG_DQ_TXDATA_OUT_net_0[151:151];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT152to152[152]       = IOG_DQ_TXDATA_OUT_net_0[152:152];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT153to153[153]       = IOG_DQ_TXDATA_OUT_net_0[153:153];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT154to154[154]       = IOG_DQ_TXDATA_OUT_net_0[154:154];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT155to155[155]       = IOG_DQ_TXDATA_OUT_net_0[155:155];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT156to156[156]       = IOG_DQ_TXDATA_OUT_net_0[156:156];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT157to157[157]       = IOG_DQ_TXDATA_OUT_net_0[157:157];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT158to158[158]       = IOG_DQ_TXDATA_OUT_net_0[158:158];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT159to159[159]       = IOG_DQ_TXDATA_OUT_net_0[159:159];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT160to160[160]       = IOG_DQ_TXDATA_OUT_net_0[160:160];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT161to161[161]       = IOG_DQ_TXDATA_OUT_net_0[161:161];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT162to162[162]       = IOG_DQ_TXDATA_OUT_net_0[162:162];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT163to163[163]       = IOG_DQ_TXDATA_OUT_net_0[163:163];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT164to164[164]       = IOG_DQ_TXDATA_OUT_net_0[164:164];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT165to165[165]       = IOG_DQ_TXDATA_OUT_net_0[165:165];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT166to166[166]       = IOG_DQ_TXDATA_OUT_net_0[166:166];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT167to167[167]       = IOG_DQ_TXDATA_OUT_net_0[167:167];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT168to168[168]       = IOG_DQ_TXDATA_OUT_net_0[168:168];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT169to169[169]       = IOG_DQ_TXDATA_OUT_net_0[169:169];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT170to170[170]       = IOG_DQ_TXDATA_OUT_net_0[170:170];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT171to171[171]       = IOG_DQ_TXDATA_OUT_net_0[171:171];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT172to172[172]       = IOG_DQ_TXDATA_OUT_net_0[172:172];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT173to173[173]       = IOG_DQ_TXDATA_OUT_net_0[173:173];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT174to174[174]       = IOG_DQ_TXDATA_OUT_net_0[174:174];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT175to175[175]       = IOG_DQ_TXDATA_OUT_net_0[175:175];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT176to176[176]       = IOG_DQ_TXDATA_OUT_net_0[176:176];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT177to177[177]       = IOG_DQ_TXDATA_OUT_net_0[177:177];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT178to178[178]       = IOG_DQ_TXDATA_OUT_net_0[178:178];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT179to179[179]       = IOG_DQ_TXDATA_OUT_net_0[179:179];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT180to180[180]       = IOG_DQ_TXDATA_OUT_net_0[180:180];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT181to181[181]       = IOG_DQ_TXDATA_OUT_net_0[181:181];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT182to182[182]       = IOG_DQ_TXDATA_OUT_net_0[182:182];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT183to183[183]       = IOG_DQ_TXDATA_OUT_net_0[183:183];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT184to184[184]       = IOG_DQ_TXDATA_OUT_net_0[184:184];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT185to185[185]       = IOG_DQ_TXDATA_OUT_net_0[185:185];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT186to186[186]       = IOG_DQ_TXDATA_OUT_net_0[186:186];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT187to187[187]       = IOG_DQ_TXDATA_OUT_net_0[187:187];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT188to188[188]       = IOG_DQ_TXDATA_OUT_net_0[188:188];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT189to189[189]       = IOG_DQ_TXDATA_OUT_net_0[189:189];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT190to190[190]       = IOG_DQ_TXDATA_OUT_net_0[190:190];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT191to191[191]       = IOG_DQ_TXDATA_OUT_net_0[191:191];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT192to192[192]       = IOG_DQ_TXDATA_OUT_net_0[192:192];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT193to193[193]       = IOG_DQ_TXDATA_OUT_net_0[193:193];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT194to194[194]       = IOG_DQ_TXDATA_OUT_net_0[194:194];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT195to195[195]       = IOG_DQ_TXDATA_OUT_net_0[195:195];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT196to196[196]       = IOG_DQ_TXDATA_OUT_net_0[196:196];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT197to197[197]       = IOG_DQ_TXDATA_OUT_net_0[197:197];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT198to198[198]       = IOG_DQ_TXDATA_OUT_net_0[198:198];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT199to199[199]       = IOG_DQ_TXDATA_OUT_net_0[199:199];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT200to200[200]       = IOG_DQ_TXDATA_OUT_net_0[200:200];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT201to201[201]       = IOG_DQ_TXDATA_OUT_net_0[201:201];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT202to202[202]       = IOG_DQ_TXDATA_OUT_net_0[202:202];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT203to203[203]       = IOG_DQ_TXDATA_OUT_net_0[203:203];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT204to204[204]       = IOG_DQ_TXDATA_OUT_net_0[204:204];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT205to205[205]       = IOG_DQ_TXDATA_OUT_net_0[205:205];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT206to206[206]       = IOG_DQ_TXDATA_OUT_net_0[206:206];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT207to207[207]       = IOG_DQ_TXDATA_OUT_net_0[207:207];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT208to208[208]       = IOG_DQ_TXDATA_OUT_net_0[208:208];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT209to209[209]       = IOG_DQ_TXDATA_OUT_net_0[209:209];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT210to210[210]       = IOG_DQ_TXDATA_OUT_net_0[210:210];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT211to211[211]       = IOG_DQ_TXDATA_OUT_net_0[211:211];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT212to212[212]       = IOG_DQ_TXDATA_OUT_net_0[212:212];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT213to213[213]       = IOG_DQ_TXDATA_OUT_net_0[213:213];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT214to214[214]       = IOG_DQ_TXDATA_OUT_net_0[214:214];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT215to215[215]       = IOG_DQ_TXDATA_OUT_net_0[215:215];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT216to216[216]       = IOG_DQ_TXDATA_OUT_net_0[216:216];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT217to217[217]       = IOG_DQ_TXDATA_OUT_net_0[217:217];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT218to218[218]       = IOG_DQ_TXDATA_OUT_net_0[218:218];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT219to219[219]       = IOG_DQ_TXDATA_OUT_net_0[219:219];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT220to220[220]       = IOG_DQ_TXDATA_OUT_net_0[220:220];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT221to221[221]       = IOG_DQ_TXDATA_OUT_net_0[221:221];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT222to222[222]       = IOG_DQ_TXDATA_OUT_net_0[222:222];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT223to223[223]       = IOG_DQ_TXDATA_OUT_net_0[223:223];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT224to224[224]       = IOG_DQ_TXDATA_OUT_net_0[224:224];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT225to225[225]       = IOG_DQ_TXDATA_OUT_net_0[225:225];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT226to226[226]       = IOG_DQ_TXDATA_OUT_net_0[226:226];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT227to227[227]       = IOG_DQ_TXDATA_OUT_net_0[227:227];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT228to228[228]       = IOG_DQ_TXDATA_OUT_net_0[228:228];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT229to229[229]       = IOG_DQ_TXDATA_OUT_net_0[229:229];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT230to230[230]       = IOG_DQ_TXDATA_OUT_net_0[230:230];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT231to231[231]       = IOG_DQ_TXDATA_OUT_net_0[231:231];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT232to232[232]       = IOG_DQ_TXDATA_OUT_net_0[232:232];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT233to233[233]       = IOG_DQ_TXDATA_OUT_net_0[233:233];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT234to234[234]       = IOG_DQ_TXDATA_OUT_net_0[234:234];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT235to235[235]       = IOG_DQ_TXDATA_OUT_net_0[235:235];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT236to236[236]       = IOG_DQ_TXDATA_OUT_net_0[236:236];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT237to237[237]       = IOG_DQ_TXDATA_OUT_net_0[237:237];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT238to238[238]       = IOG_DQ_TXDATA_OUT_net_0[238:238];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT239to239[239]       = IOG_DQ_TXDATA_OUT_net_0[239:239];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT240to240[240]       = IOG_DQ_TXDATA_OUT_net_0[240:240];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT241to241[241]       = IOG_DQ_TXDATA_OUT_net_0[241:241];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT242to242[242]       = IOG_DQ_TXDATA_OUT_net_0[242:242];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT243to243[243]       = IOG_DQ_TXDATA_OUT_net_0[243:243];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT244to244[244]       = IOG_DQ_TXDATA_OUT_net_0[244:244];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT245to245[245]       = IOG_DQ_TXDATA_OUT_net_0[245:245];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT246to246[246]       = IOG_DQ_TXDATA_OUT_net_0[246:246];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT247to247[247]       = IOG_DQ_TXDATA_OUT_net_0[247:247];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT248to248[248]       = IOG_DQ_TXDATA_OUT_net_0[248:248];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT249to249[249]       = IOG_DQ_TXDATA_OUT_net_0[249:249];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT250to250[250]       = IOG_DQ_TXDATA_OUT_net_0[250:250];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT251to251[251]       = IOG_DQ_TXDATA_OUT_net_0[251:251];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT252to252[252]       = IOG_DQ_TXDATA_OUT_net_0[252:252];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT253to253[253]       = IOG_DQ_TXDATA_OUT_net_0[253:253];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT254to254[254]       = IOG_DQ_TXDATA_OUT_net_0[254:254];
assign IOD_TRAINING_0_IOG_DQ_TXDATA_OUT255to255[255]       = IOG_DQ_TXDATA_OUT_net_0[255:255];
assign IOD_TRAINING_0_IOG_OE_P00to0[0]                     = IOG_OE_P0_net_0[0:0];
assign IOD_TRAINING_0_IOG_OE_P01to1[1]                     = IOG_OE_P0_net_0[1:1];
assign IOD_TRAINING_0_IOG_OE_P02to2[2]                     = IOG_OE_P0_net_0[2:2];
assign IOD_TRAINING_0_IOG_OE_P03to3[3]                     = IOG_OE_P0_net_0[3:3];
assign IOD_TRAINING_0_IOG_OE_P10to0[0]                     = IOG_OE_P1_net_0[0:0];
assign IOD_TRAINING_0_IOG_OE_P11to1[1]                     = IOG_OE_P1_net_0[1:1];
assign IOD_TRAINING_0_IOG_OE_P12to2[2]                     = IOG_OE_P1_net_0[2:2];
assign IOD_TRAINING_0_IOG_OE_P13to3[3]                     = IOG_OE_P1_net_0[3:3];
assign IOD_TRAINING_0_IOG_OE_P20to0[0]                     = IOG_OE_P2_net_0[0:0];
assign IOD_TRAINING_0_IOG_OE_P21to1[1]                     = IOG_OE_P2_net_0[1:1];
assign IOD_TRAINING_0_IOG_OE_P22to2[2]                     = IOG_OE_P2_net_0[2:2];
assign IOD_TRAINING_0_IOG_OE_P23to3[3]                     = IOG_OE_P2_net_0[3:3];
assign IOD_TRAINING_0_IOG_OE_P30to0[0]                     = IOG_OE_P3_net_0[0:0];
assign IOD_TRAINING_0_IOG_OE_P31to1[1]                     = IOG_OE_P3_net_0[1:1];
assign IOD_TRAINING_0_IOG_OE_P32to2[2]                     = IOG_OE_P3_net_0[2:2];
assign IOD_TRAINING_0_IOG_OE_P33to3[3]                     = IOG_OE_P3_net_0[3:3];
assign IOD_TRAINING_0_IOG_RDDATA_EN_P0_N0to0[0]            = IOG_RDDATA_EN_P0_N_net_0[0:0];
assign IOD_TRAINING_0_IOG_RDDATA_EN_P0_N1to1[1]            = IOG_RDDATA_EN_P0_N_net_0[1:1];
assign IOD_TRAINING_0_IOG_RDDATA_EN_P0_N2to2[2]            = IOG_RDDATA_EN_P0_N_net_0[2:2];
assign IOD_TRAINING_0_IOG_RDDATA_EN_P0_N3to3[3]            = IOG_RDDATA_EN_P0_N_net_0[3:3];
assign IOD_TRAINING_0_IOG_RDDATA_EN_P0_P0to0[0]            = IOG_RDDATA_EN_P0_P_net_0[0:0];
assign IOD_TRAINING_0_IOG_RDDATA_EN_P0_P1to1[1]            = IOG_RDDATA_EN_P0_P_net_0[1:1];
assign IOD_TRAINING_0_IOG_RDDATA_EN_P0_P2to2[2]            = IOG_RDDATA_EN_P0_P_net_0[2:2];
assign IOD_TRAINING_0_IOG_RDDATA_EN_P0_P3to3[3]            = IOG_RDDATA_EN_P0_P_net_0[3:3];
assign IOD_TRAINING_0_IOG_RDDATA_EN_P1_N0to0[0]            = IOG_RDDATA_EN_P1_N_net_0[0:0];
assign IOD_TRAINING_0_IOG_RDDATA_EN_P1_N1to1[1]            = IOG_RDDATA_EN_P1_N_net_0[1:1];
assign IOD_TRAINING_0_IOG_RDDATA_EN_P1_N2to2[2]            = IOG_RDDATA_EN_P1_N_net_0[2:2];
assign IOD_TRAINING_0_IOG_RDDATA_EN_P1_N3to3[3]            = IOG_RDDATA_EN_P1_N_net_0[3:3];
assign IOD_TRAINING_0_IOG_RDDATA_EN_P1_P0to0[0]            = IOG_RDDATA_EN_P1_P_net_0[0:0];
assign IOD_TRAINING_0_IOG_RDDATA_EN_P1_P1to1[1]            = IOG_RDDATA_EN_P1_P_net_0[1:1];
assign IOD_TRAINING_0_IOG_RDDATA_EN_P1_P2to2[2]            = IOG_RDDATA_EN_P1_P_net_0[2:2];
assign IOD_TRAINING_0_IOG_RDDATA_EN_P1_P3to3[3]            = IOG_RDDATA_EN_P1_P_net_0[3:3];
assign IOD_TRAINING_0_IOG_RDDATA_EN_P2_N0to0[0]            = IOG_RDDATA_EN_P2_N_net_0[0:0];
assign IOD_TRAINING_0_IOG_RDDATA_EN_P2_N1to1[1]            = IOG_RDDATA_EN_P2_N_net_0[1:1];
assign IOD_TRAINING_0_IOG_RDDATA_EN_P2_N2to2[2]            = IOG_RDDATA_EN_P2_N_net_0[2:2];
assign IOD_TRAINING_0_IOG_RDDATA_EN_P2_N3to3[3]            = IOG_RDDATA_EN_P2_N_net_0[3:3];
assign IOD_TRAINING_0_IOG_RDDATA_EN_P2_P0to0[0]            = IOG_RDDATA_EN_P2_P_net_0[0:0];
assign IOD_TRAINING_0_IOG_RDDATA_EN_P2_P1to1[1]            = IOG_RDDATA_EN_P2_P_net_0[1:1];
assign IOD_TRAINING_0_IOG_RDDATA_EN_P2_P2to2[2]            = IOG_RDDATA_EN_P2_P_net_0[2:2];
assign IOD_TRAINING_0_IOG_RDDATA_EN_P2_P3to3[3]            = IOG_RDDATA_EN_P2_P_net_0[3:3];
assign IOD_TRAINING_0_IOG_RDDATA_EN_P3_N0to0[0]            = IOG_RDDATA_EN_P3_N_net_0[0:0];
assign IOD_TRAINING_0_IOG_RDDATA_EN_P3_N1to1[1]            = IOG_RDDATA_EN_P3_N_net_0[1:1];
assign IOD_TRAINING_0_IOG_RDDATA_EN_P3_N2to2[2]            = IOG_RDDATA_EN_P3_N_net_0[2:2];
assign IOD_TRAINING_0_IOG_RDDATA_EN_P3_N3to3[3]            = IOG_RDDATA_EN_P3_N_net_0[3:3];
assign IOD_TRAINING_0_IOG_RDDATA_EN_P3_P0to0[0]            = IOG_RDDATA_EN_P3_P_net_0[0:0];
assign IOD_TRAINING_0_IOG_RDDATA_EN_P3_P1to1[1]            = IOG_RDDATA_EN_P3_P_net_0[1:1];
assign IOD_TRAINING_0_IOG_RDDATA_EN_P3_P2to2[2]            = IOG_RDDATA_EN_P3_P_net_0[2:2];
assign IOD_TRAINING_0_IOG_RDDATA_EN_P3_P3to3[3]            = IOG_RDDATA_EN_P3_P_net_0[3:3];
assign IOD_TRAINING_0_LOAD0to0[0]                          = LOAD_net_0[0:0];
assign IOD_TRAINING_0_LOAD1to1[1]                          = LOAD_net_0[1:1];
assign IOD_TRAINING_0_LOAD2to2[2]                          = LOAD_net_0[2:2];
assign IOD_TRAINING_0_LOAD3to3[3]                          = LOAD_net_0[3:3];
assign IOD_TRAINING_0_LOAD4to4[4]                          = LOAD_net_0[4:4];
assign IOD_TRAINING_0_LOAD5to5[5]                          = LOAD_net_0[5:5];
assign IOD_TRAINING_0_LOAD6to6[6]                          = LOAD_net_0[6:6];
assign IOD_TRAINING_0_LOAD7to7[7]                          = LOAD_net_0[7:7];
assign IOD_TRAINING_0_LOAD8to8[8]                          = LOAD_net_0[8:8];
assign IOD_TRAINING_0_LOAD9to9[9]                          = LOAD_net_0[9:9];
assign IOD_TRAINING_0_LOAD10to10[10]                       = LOAD_net_0[10:10];
assign IOD_TRAINING_0_LOAD11to11[11]                       = LOAD_net_0[11:11];
assign IOD_TRAINING_0_LOAD12to12[12]                       = LOAD_net_0[12:12];
assign IOD_TRAINING_0_LOAD13to13[13]                       = LOAD_net_0[13:13];
assign IOD_TRAINING_0_LOAD14to14[14]                       = LOAD_net_0[14:14];
assign IOD_TRAINING_0_LOAD15to15[15]                       = LOAD_net_0[15:15];
assign IOD_TRAINING_0_LOAD16to16[16]                       = LOAD_net_0[16:16];
assign IOD_TRAINING_0_LOAD17to17[17]                       = LOAD_net_0[17:17];
assign IOD_TRAINING_0_LOAD18to18[18]                       = LOAD_net_0[18:18];
assign IOD_TRAINING_0_LOAD19to19[19]                       = LOAD_net_0[19:19];
assign IOD_TRAINING_0_LOAD20to20[20]                       = LOAD_net_0[20:20];
assign IOD_TRAINING_0_LOAD21to21[21]                       = LOAD_net_0[21:21];
assign IOD_TRAINING_0_LOAD22to22[22]                       = LOAD_net_0[22:22];
assign IOD_TRAINING_0_LOAD23to23[23]                       = LOAD_net_0[23:23];
assign IOD_TRAINING_0_LOAD24to24[24]                       = LOAD_net_0[24:24];
assign IOD_TRAINING_0_LOAD25to25[25]                       = LOAD_net_0[25:25];
assign IOD_TRAINING_0_LOAD26to26[26]                       = LOAD_net_0[26:26];
assign IOD_TRAINING_0_LOAD27to27[27]                       = LOAD_net_0[27:27];
assign IOD_TRAINING_0_LOAD28to28[28]                       = LOAD_net_0[28:28];
assign IOD_TRAINING_0_LOAD29to29[29]                       = LOAD_net_0[29:29];
assign IOD_TRAINING_0_LOAD30to30[30]                       = LOAD_net_0[30:30];
assign IOD_TRAINING_0_LOAD31to31[31]                       = LOAD_net_0[31:31];
assign IOD_TRAINING_0_LOAD32to32[32]                       = LOAD_net_0[32:32];
assign IOD_TRAINING_0_LOAD33to33[33]                       = LOAD_net_0[33:33];
assign IOD_TRAINING_0_LOAD34to34[34]                       = LOAD_net_0[34:34];
assign IOD_TRAINING_0_LOAD35to35[35]                       = LOAD_net_0[35:35];
assign IOD_TRAINING_0_MOVE0to0[0]                          = MOVE_net_0[0:0];
assign IOD_TRAINING_0_MOVE1to1[1]                          = MOVE_net_0[1:1];
assign IOD_TRAINING_0_MOVE2to2[2]                          = MOVE_net_0[2:2];
assign IOD_TRAINING_0_MOVE3to3[3]                          = MOVE_net_0[3:3];
assign IOD_TRAINING_0_MOVE4to4[4]                          = MOVE_net_0[4:4];
assign IOD_TRAINING_0_MOVE5to5[5]                          = MOVE_net_0[5:5];
assign IOD_TRAINING_0_MOVE6to6[6]                          = MOVE_net_0[6:6];
assign IOD_TRAINING_0_MOVE7to7[7]                          = MOVE_net_0[7:7];
assign IOD_TRAINING_0_MOVE8to8[8]                          = MOVE_net_0[8:8];
assign IOD_TRAINING_0_MOVE9to9[9]                          = MOVE_net_0[9:9];
assign IOD_TRAINING_0_MOVE10to10[10]                       = MOVE_net_0[10:10];
assign IOD_TRAINING_0_MOVE11to11[11]                       = MOVE_net_0[11:11];
assign IOD_TRAINING_0_MOVE12to12[12]                       = MOVE_net_0[12:12];
assign IOD_TRAINING_0_MOVE13to13[13]                       = MOVE_net_0[13:13];
assign IOD_TRAINING_0_MOVE14to14[14]                       = MOVE_net_0[14:14];
assign IOD_TRAINING_0_MOVE15to15[15]                       = MOVE_net_0[15:15];
assign IOD_TRAINING_0_MOVE16to16[16]                       = MOVE_net_0[16:16];
assign IOD_TRAINING_0_MOVE17to17[17]                       = MOVE_net_0[17:17];
assign IOD_TRAINING_0_MOVE18to18[18]                       = MOVE_net_0[18:18];
assign IOD_TRAINING_0_MOVE19to19[19]                       = MOVE_net_0[19:19];
assign IOD_TRAINING_0_MOVE20to20[20]                       = MOVE_net_0[20:20];
assign IOD_TRAINING_0_MOVE21to21[21]                       = MOVE_net_0[21:21];
assign IOD_TRAINING_0_MOVE22to22[22]                       = MOVE_net_0[22:22];
assign IOD_TRAINING_0_MOVE23to23[23]                       = MOVE_net_0[23:23];
assign IOD_TRAINING_0_MOVE24to24[24]                       = MOVE_net_0[24:24];
assign IOD_TRAINING_0_MOVE25to25[25]                       = MOVE_net_0[25:25];
assign IOD_TRAINING_0_MOVE26to26[26]                       = MOVE_net_0[26:26];
assign IOD_TRAINING_0_MOVE27to27[27]                       = MOVE_net_0[27:27];
assign IOD_TRAINING_0_MOVE28to28[28]                       = MOVE_net_0[28:28];
assign IOD_TRAINING_0_MOVE29to29[29]                       = MOVE_net_0[29:29];
assign IOD_TRAINING_0_MOVE30to30[30]                       = MOVE_net_0[30:30];
assign IOD_TRAINING_0_MOVE31to31[31]                       = MOVE_net_0[31:31];
assign IOD_TRAINING_0_MOVE32to32[32]                       = MOVE_net_0[32:32];
assign IOD_TRAINING_0_MOVE33to33[33]                       = MOVE_net_0[33:33];
assign IOD_TRAINING_0_MOVE34to34[34]                       = MOVE_net_0[34:34];
assign IOD_TRAINING_0_MOVE35to35[35]                       = MOVE_net_0[35:35];
assign LANE_0_IOD_DQ_RX_DATA_00to0[0]                      = RX_DATA_0_net_3[0:0];
assign LANE_0_IOD_DQ_RX_DATA_01to1[1]                      = RX_DATA_0_net_3[1:1];
assign LANE_0_IOD_DQ_RX_DATA_02to2[2]                      = RX_DATA_0_net_3[2:2];
assign LANE_0_IOD_DQ_RX_DATA_03to3[3]                      = RX_DATA_0_net_3[3:3];
assign LANE_0_IOD_DQ_RX_DATA_04to4[4]                      = RX_DATA_0_net_3[4:4];
assign LANE_0_IOD_DQ_RX_DATA_05to5[5]                      = RX_DATA_0_net_3[5:5];
assign LANE_0_IOD_DQ_RX_DATA_06to6[6]                      = RX_DATA_0_net_3[6:6];
assign LANE_0_IOD_DQ_RX_DATA_07to7[7]                      = RX_DATA_0_net_3[7:7];
assign LANE_0_IOD_DQ_RX_DATA_10to0[0]                      = RX_DATA_1_net_0[0:0];
assign LANE_0_IOD_DQ_RX_DATA_11to1[1]                      = RX_DATA_1_net_0[1:1];
assign LANE_0_IOD_DQ_RX_DATA_12to2[2]                      = RX_DATA_1_net_0[2:2];
assign LANE_0_IOD_DQ_RX_DATA_13to3[3]                      = RX_DATA_1_net_0[3:3];
assign LANE_0_IOD_DQ_RX_DATA_14to4[4]                      = RX_DATA_1_net_0[4:4];
assign LANE_0_IOD_DQ_RX_DATA_15to5[5]                      = RX_DATA_1_net_0[5:5];
assign LANE_0_IOD_DQ_RX_DATA_16to6[6]                      = RX_DATA_1_net_0[6:6];
assign LANE_0_IOD_DQ_RX_DATA_17to7[7]                      = RX_DATA_1_net_0[7:7];
assign LANE_0_IOD_DQ_RX_DATA_20to0[0]                      = RX_DATA_2_net_0[0:0];
assign LANE_0_IOD_DQ_RX_DATA_21to1[1]                      = RX_DATA_2_net_0[1:1];
assign LANE_0_IOD_DQ_RX_DATA_22to2[2]                      = RX_DATA_2_net_0[2:2];
assign LANE_0_IOD_DQ_RX_DATA_23to3[3]                      = RX_DATA_2_net_0[3:3];
assign LANE_0_IOD_DQ_RX_DATA_24to4[4]                      = RX_DATA_2_net_0[4:4];
assign LANE_0_IOD_DQ_RX_DATA_25to5[5]                      = RX_DATA_2_net_0[5:5];
assign LANE_0_IOD_DQ_RX_DATA_26to6[6]                      = RX_DATA_2_net_0[6:6];
assign LANE_0_IOD_DQ_RX_DATA_27to7[7]                      = RX_DATA_2_net_0[7:7];
assign LANE_0_IOD_DQ_RX_DATA_30to0[0]                      = RX_DATA_3_net_0[0:0];
assign LANE_0_IOD_DQ_RX_DATA_31to1[1]                      = RX_DATA_3_net_0[1:1];
assign LANE_0_IOD_DQ_RX_DATA_32to2[2]                      = RX_DATA_3_net_0[2:2];
assign LANE_0_IOD_DQ_RX_DATA_33to3[3]                      = RX_DATA_3_net_0[3:3];
assign LANE_0_IOD_DQ_RX_DATA_34to4[4]                      = RX_DATA_3_net_0[4:4];
assign LANE_0_IOD_DQ_RX_DATA_35to5[5]                      = RX_DATA_3_net_0[5:5];
assign LANE_0_IOD_DQ_RX_DATA_36to6[6]                      = RX_DATA_3_net_0[6:6];
assign LANE_0_IOD_DQ_RX_DATA_37to7[7]                      = RX_DATA_3_net_0[7:7];
assign LANE_0_IOD_DQ_RX_DATA_40to0[0]                      = RX_DATA_4_net_0[0:0];
assign LANE_0_IOD_DQ_RX_DATA_41to1[1]                      = RX_DATA_4_net_0[1:1];
assign LANE_0_IOD_DQ_RX_DATA_42to2[2]                      = RX_DATA_4_net_0[2:2];
assign LANE_0_IOD_DQ_RX_DATA_43to3[3]                      = RX_DATA_4_net_0[3:3];
assign LANE_0_IOD_DQ_RX_DATA_44to4[4]                      = RX_DATA_4_net_0[4:4];
assign LANE_0_IOD_DQ_RX_DATA_45to5[5]                      = RX_DATA_4_net_0[5:5];
assign LANE_0_IOD_DQ_RX_DATA_46to6[6]                      = RX_DATA_4_net_0[6:6];
assign LANE_0_IOD_DQ_RX_DATA_47to7[7]                      = RX_DATA_4_net_0[7:7];
assign LANE_0_IOD_DQ_RX_DATA_50to0[0]                      = RX_DATA_5_net_0[0:0];
assign LANE_0_IOD_DQ_RX_DATA_51to1[1]                      = RX_DATA_5_net_0[1:1];
assign LANE_0_IOD_DQ_RX_DATA_52to2[2]                      = RX_DATA_5_net_0[2:2];
assign LANE_0_IOD_DQ_RX_DATA_53to3[3]                      = RX_DATA_5_net_0[3:3];
assign LANE_0_IOD_DQ_RX_DATA_54to4[4]                      = RX_DATA_5_net_0[4:4];
assign LANE_0_IOD_DQ_RX_DATA_55to5[5]                      = RX_DATA_5_net_0[5:5];
assign LANE_0_IOD_DQ_RX_DATA_56to6[6]                      = RX_DATA_5_net_0[6:6];
assign LANE_0_IOD_DQ_RX_DATA_57to7[7]                      = RX_DATA_5_net_0[7:7];
assign LANE_0_IOD_DQ_RX_DATA_60to0[0]                      = RX_DATA_6_net_0[0:0];
assign LANE_0_IOD_DQ_RX_DATA_61to1[1]                      = RX_DATA_6_net_0[1:1];
assign LANE_0_IOD_DQ_RX_DATA_62to2[2]                      = RX_DATA_6_net_0[2:2];
assign LANE_0_IOD_DQ_RX_DATA_63to3[3]                      = RX_DATA_6_net_0[3:3];
assign LANE_0_IOD_DQ_RX_DATA_64to4[4]                      = RX_DATA_6_net_0[4:4];
assign LANE_0_IOD_DQ_RX_DATA_65to5[5]                      = RX_DATA_6_net_0[5:5];
assign LANE_0_IOD_DQ_RX_DATA_66to6[6]                      = RX_DATA_6_net_0[6:6];
assign LANE_0_IOD_DQ_RX_DATA_67to7[7]                      = RX_DATA_6_net_0[7:7];
assign LANE_0_IOD_DQ_RX_DATA_70to0[0]                      = RX_DATA_7_net_0[0:0];
assign LANE_0_IOD_DQ_RX_DATA_71to1[1]                      = RX_DATA_7_net_0[1:1];
assign LANE_0_IOD_DQ_RX_DATA_72to2[2]                      = RX_DATA_7_net_0[2:2];
assign LANE_0_IOD_DQ_RX_DATA_73to3[3]                      = RX_DATA_7_net_0[3:3];
assign LANE_0_IOD_DQ_RX_DATA_74to4[4]                      = RX_DATA_7_net_0[4:4];
assign LANE_0_IOD_DQ_RX_DATA_75to5[5]                      = RX_DATA_7_net_0[5:5];
assign LANE_0_IOD_DQ_RX_DATA_76to6[6]                      = RX_DATA_7_net_0[6:6];
assign LANE_0_IOD_DQ_RX_DATA_77to7[7]                      = RX_DATA_7_net_0[7:7];
assign LANE_0_IOD_DQSW_TRAINING_RX_DATA_00to0[0]           = RX_DATA_0_net_4[0:0];
assign LANE_0_IOD_DQSW_TRAINING_RX_DATA_01to1[1]           = RX_DATA_0_net_4[1:1];
assign LANE_0_IOD_READ_TRAINING_RX_DATA_06to6[6]           = RX_DATA_0_net_5[6:6];
assign LANE_0_IOD_READ_TRAINING_RX_DATA_07to7[7]           = RX_DATA_0_net_5[7:7];
assign LANE_1_IOD_DQ_RX_DATA_00to0[0]                      = RX_DATA_0_net_6[0:0];
assign LANE_1_IOD_DQ_RX_DATA_01to1[1]                      = RX_DATA_0_net_6[1:1];
assign LANE_1_IOD_DQ_RX_DATA_02to2[2]                      = RX_DATA_0_net_6[2:2];
assign LANE_1_IOD_DQ_RX_DATA_03to3[3]                      = RX_DATA_0_net_6[3:3];
assign LANE_1_IOD_DQ_RX_DATA_04to4[4]                      = RX_DATA_0_net_6[4:4];
assign LANE_1_IOD_DQ_RX_DATA_05to5[5]                      = RX_DATA_0_net_6[5:5];
assign LANE_1_IOD_DQ_RX_DATA_06to6[6]                      = RX_DATA_0_net_6[6:6];
assign LANE_1_IOD_DQ_RX_DATA_07to7[7]                      = RX_DATA_0_net_6[7:7];
assign LANE_1_IOD_DQ_RX_DATA_10to0[0]                      = RX_DATA_1_net_1[0:0];
assign LANE_1_IOD_DQ_RX_DATA_11to1[1]                      = RX_DATA_1_net_1[1:1];
assign LANE_1_IOD_DQ_RX_DATA_12to2[2]                      = RX_DATA_1_net_1[2:2];
assign LANE_1_IOD_DQ_RX_DATA_13to3[3]                      = RX_DATA_1_net_1[3:3];
assign LANE_1_IOD_DQ_RX_DATA_14to4[4]                      = RX_DATA_1_net_1[4:4];
assign LANE_1_IOD_DQ_RX_DATA_15to5[5]                      = RX_DATA_1_net_1[5:5];
assign LANE_1_IOD_DQ_RX_DATA_16to6[6]                      = RX_DATA_1_net_1[6:6];
assign LANE_1_IOD_DQ_RX_DATA_17to7[7]                      = RX_DATA_1_net_1[7:7];
assign LANE_1_IOD_DQ_RX_DATA_20to0[0]                      = RX_DATA_2_net_1[0:0];
assign LANE_1_IOD_DQ_RX_DATA_21to1[1]                      = RX_DATA_2_net_1[1:1];
assign LANE_1_IOD_DQ_RX_DATA_22to2[2]                      = RX_DATA_2_net_1[2:2];
assign LANE_1_IOD_DQ_RX_DATA_23to3[3]                      = RX_DATA_2_net_1[3:3];
assign LANE_1_IOD_DQ_RX_DATA_24to4[4]                      = RX_DATA_2_net_1[4:4];
assign LANE_1_IOD_DQ_RX_DATA_25to5[5]                      = RX_DATA_2_net_1[5:5];
assign LANE_1_IOD_DQ_RX_DATA_26to6[6]                      = RX_DATA_2_net_1[6:6];
assign LANE_1_IOD_DQ_RX_DATA_27to7[7]                      = RX_DATA_2_net_1[7:7];
assign LANE_1_IOD_DQ_RX_DATA_30to0[0]                      = RX_DATA_3_net_1[0:0];
assign LANE_1_IOD_DQ_RX_DATA_31to1[1]                      = RX_DATA_3_net_1[1:1];
assign LANE_1_IOD_DQ_RX_DATA_32to2[2]                      = RX_DATA_3_net_1[2:2];
assign LANE_1_IOD_DQ_RX_DATA_33to3[3]                      = RX_DATA_3_net_1[3:3];
assign LANE_1_IOD_DQ_RX_DATA_34to4[4]                      = RX_DATA_3_net_1[4:4];
assign LANE_1_IOD_DQ_RX_DATA_35to5[5]                      = RX_DATA_3_net_1[5:5];
assign LANE_1_IOD_DQ_RX_DATA_36to6[6]                      = RX_DATA_3_net_1[6:6];
assign LANE_1_IOD_DQ_RX_DATA_37to7[7]                      = RX_DATA_3_net_1[7:7];
assign LANE_1_IOD_DQ_RX_DATA_40to0[0]                      = RX_DATA_4_net_1[0:0];
assign LANE_1_IOD_DQ_RX_DATA_41to1[1]                      = RX_DATA_4_net_1[1:1];
assign LANE_1_IOD_DQ_RX_DATA_42to2[2]                      = RX_DATA_4_net_1[2:2];
assign LANE_1_IOD_DQ_RX_DATA_43to3[3]                      = RX_DATA_4_net_1[3:3];
assign LANE_1_IOD_DQ_RX_DATA_44to4[4]                      = RX_DATA_4_net_1[4:4];
assign LANE_1_IOD_DQ_RX_DATA_45to5[5]                      = RX_DATA_4_net_1[5:5];
assign LANE_1_IOD_DQ_RX_DATA_46to6[6]                      = RX_DATA_4_net_1[6:6];
assign LANE_1_IOD_DQ_RX_DATA_47to7[7]                      = RX_DATA_4_net_1[7:7];
assign LANE_1_IOD_DQ_RX_DATA_50to0[0]                      = RX_DATA_5_net_1[0:0];
assign LANE_1_IOD_DQ_RX_DATA_51to1[1]                      = RX_DATA_5_net_1[1:1];
assign LANE_1_IOD_DQ_RX_DATA_52to2[2]                      = RX_DATA_5_net_1[2:2];
assign LANE_1_IOD_DQ_RX_DATA_53to3[3]                      = RX_DATA_5_net_1[3:3];
assign LANE_1_IOD_DQ_RX_DATA_54to4[4]                      = RX_DATA_5_net_1[4:4];
assign LANE_1_IOD_DQ_RX_DATA_55to5[5]                      = RX_DATA_5_net_1[5:5];
assign LANE_1_IOD_DQ_RX_DATA_56to6[6]                      = RX_DATA_5_net_1[6:6];
assign LANE_1_IOD_DQ_RX_DATA_57to7[7]                      = RX_DATA_5_net_1[7:7];
assign LANE_1_IOD_DQ_RX_DATA_60to0[0]                      = RX_DATA_6_net_1[0:0];
assign LANE_1_IOD_DQ_RX_DATA_61to1[1]                      = RX_DATA_6_net_1[1:1];
assign LANE_1_IOD_DQ_RX_DATA_62to2[2]                      = RX_DATA_6_net_1[2:2];
assign LANE_1_IOD_DQ_RX_DATA_63to3[3]                      = RX_DATA_6_net_1[3:3];
assign LANE_1_IOD_DQ_RX_DATA_64to4[4]                      = RX_DATA_6_net_1[4:4];
assign LANE_1_IOD_DQ_RX_DATA_65to5[5]                      = RX_DATA_6_net_1[5:5];
assign LANE_1_IOD_DQ_RX_DATA_66to6[6]                      = RX_DATA_6_net_1[6:6];
assign LANE_1_IOD_DQ_RX_DATA_67to7[7]                      = RX_DATA_6_net_1[7:7];
assign LANE_1_IOD_DQ_RX_DATA_70to0[0]                      = RX_DATA_7_net_1[0:0];
assign LANE_1_IOD_DQ_RX_DATA_71to1[1]                      = RX_DATA_7_net_1[1:1];
assign LANE_1_IOD_DQ_RX_DATA_72to2[2]                      = RX_DATA_7_net_1[2:2];
assign LANE_1_IOD_DQ_RX_DATA_73to3[3]                      = RX_DATA_7_net_1[3:3];
assign LANE_1_IOD_DQ_RX_DATA_74to4[4]                      = RX_DATA_7_net_1[4:4];
assign LANE_1_IOD_DQ_RX_DATA_75to5[5]                      = RX_DATA_7_net_1[5:5];
assign LANE_1_IOD_DQ_RX_DATA_76to6[6]                      = RX_DATA_7_net_1[6:6];
assign LANE_1_IOD_DQ_RX_DATA_77to7[7]                      = RX_DATA_7_net_1[7:7];
assign LANE_1_IOD_DQSW_TRAINING_RX_DATA_00to0[0]           = RX_DATA_0_net_7[0:0];
assign LANE_1_IOD_DQSW_TRAINING_RX_DATA_01to1[1]           = RX_DATA_0_net_7[1:1];
assign LANE_1_IOD_READ_TRAINING_RX_DATA_06to6[6]           = RX_DATA_0_net_8[6:6];
assign LANE_1_IOD_READ_TRAINING_RX_DATA_07to7[7]           = RX_DATA_0_net_8[7:7];
assign LANE_2_IOD_DQ_RX_DATA_00to0[0]                      = RX_DATA_0_net_9[0:0];
assign LANE_2_IOD_DQ_RX_DATA_01to1[1]                      = RX_DATA_0_net_9[1:1];
assign LANE_2_IOD_DQ_RX_DATA_02to2[2]                      = RX_DATA_0_net_9[2:2];
assign LANE_2_IOD_DQ_RX_DATA_03to3[3]                      = RX_DATA_0_net_9[3:3];
assign LANE_2_IOD_DQ_RX_DATA_04to4[4]                      = RX_DATA_0_net_9[4:4];
assign LANE_2_IOD_DQ_RX_DATA_05to5[5]                      = RX_DATA_0_net_9[5:5];
assign LANE_2_IOD_DQ_RX_DATA_06to6[6]                      = RX_DATA_0_net_9[6:6];
assign LANE_2_IOD_DQ_RX_DATA_07to7[7]                      = RX_DATA_0_net_9[7:7];
assign LANE_2_IOD_DQ_RX_DATA_10to0[0]                      = RX_DATA_1_net_2[0:0];
assign LANE_2_IOD_DQ_RX_DATA_11to1[1]                      = RX_DATA_1_net_2[1:1];
assign LANE_2_IOD_DQ_RX_DATA_12to2[2]                      = RX_DATA_1_net_2[2:2];
assign LANE_2_IOD_DQ_RX_DATA_13to3[3]                      = RX_DATA_1_net_2[3:3];
assign LANE_2_IOD_DQ_RX_DATA_14to4[4]                      = RX_DATA_1_net_2[4:4];
assign LANE_2_IOD_DQ_RX_DATA_15to5[5]                      = RX_DATA_1_net_2[5:5];
assign LANE_2_IOD_DQ_RX_DATA_16to6[6]                      = RX_DATA_1_net_2[6:6];
assign LANE_2_IOD_DQ_RX_DATA_17to7[7]                      = RX_DATA_1_net_2[7:7];
assign LANE_2_IOD_DQ_RX_DATA_20to0[0]                      = RX_DATA_2_net_2[0:0];
assign LANE_2_IOD_DQ_RX_DATA_21to1[1]                      = RX_DATA_2_net_2[1:1];
assign LANE_2_IOD_DQ_RX_DATA_22to2[2]                      = RX_DATA_2_net_2[2:2];
assign LANE_2_IOD_DQ_RX_DATA_23to3[3]                      = RX_DATA_2_net_2[3:3];
assign LANE_2_IOD_DQ_RX_DATA_24to4[4]                      = RX_DATA_2_net_2[4:4];
assign LANE_2_IOD_DQ_RX_DATA_25to5[5]                      = RX_DATA_2_net_2[5:5];
assign LANE_2_IOD_DQ_RX_DATA_26to6[6]                      = RX_DATA_2_net_2[6:6];
assign LANE_2_IOD_DQ_RX_DATA_27to7[7]                      = RX_DATA_2_net_2[7:7];
assign LANE_2_IOD_DQ_RX_DATA_30to0[0]                      = RX_DATA_3_net_2[0:0];
assign LANE_2_IOD_DQ_RX_DATA_31to1[1]                      = RX_DATA_3_net_2[1:1];
assign LANE_2_IOD_DQ_RX_DATA_32to2[2]                      = RX_DATA_3_net_2[2:2];
assign LANE_2_IOD_DQ_RX_DATA_33to3[3]                      = RX_DATA_3_net_2[3:3];
assign LANE_2_IOD_DQ_RX_DATA_34to4[4]                      = RX_DATA_3_net_2[4:4];
assign LANE_2_IOD_DQ_RX_DATA_35to5[5]                      = RX_DATA_3_net_2[5:5];
assign LANE_2_IOD_DQ_RX_DATA_36to6[6]                      = RX_DATA_3_net_2[6:6];
assign LANE_2_IOD_DQ_RX_DATA_37to7[7]                      = RX_DATA_3_net_2[7:7];
assign LANE_2_IOD_DQ_RX_DATA_40to0[0]                      = RX_DATA_4_net_2[0:0];
assign LANE_2_IOD_DQ_RX_DATA_41to1[1]                      = RX_DATA_4_net_2[1:1];
assign LANE_2_IOD_DQ_RX_DATA_42to2[2]                      = RX_DATA_4_net_2[2:2];
assign LANE_2_IOD_DQ_RX_DATA_43to3[3]                      = RX_DATA_4_net_2[3:3];
assign LANE_2_IOD_DQ_RX_DATA_44to4[4]                      = RX_DATA_4_net_2[4:4];
assign LANE_2_IOD_DQ_RX_DATA_45to5[5]                      = RX_DATA_4_net_2[5:5];
assign LANE_2_IOD_DQ_RX_DATA_46to6[6]                      = RX_DATA_4_net_2[6:6];
assign LANE_2_IOD_DQ_RX_DATA_47to7[7]                      = RX_DATA_4_net_2[7:7];
assign LANE_2_IOD_DQ_RX_DATA_50to0[0]                      = RX_DATA_5_net_2[0:0];
assign LANE_2_IOD_DQ_RX_DATA_51to1[1]                      = RX_DATA_5_net_2[1:1];
assign LANE_2_IOD_DQ_RX_DATA_52to2[2]                      = RX_DATA_5_net_2[2:2];
assign LANE_2_IOD_DQ_RX_DATA_53to3[3]                      = RX_DATA_5_net_2[3:3];
assign LANE_2_IOD_DQ_RX_DATA_54to4[4]                      = RX_DATA_5_net_2[4:4];
assign LANE_2_IOD_DQ_RX_DATA_55to5[5]                      = RX_DATA_5_net_2[5:5];
assign LANE_2_IOD_DQ_RX_DATA_56to6[6]                      = RX_DATA_5_net_2[6:6];
assign LANE_2_IOD_DQ_RX_DATA_57to7[7]                      = RX_DATA_5_net_2[7:7];
assign LANE_2_IOD_DQ_RX_DATA_60to0[0]                      = RX_DATA_6_net_2[0:0];
assign LANE_2_IOD_DQ_RX_DATA_61to1[1]                      = RX_DATA_6_net_2[1:1];
assign LANE_2_IOD_DQ_RX_DATA_62to2[2]                      = RX_DATA_6_net_2[2:2];
assign LANE_2_IOD_DQ_RX_DATA_63to3[3]                      = RX_DATA_6_net_2[3:3];
assign LANE_2_IOD_DQ_RX_DATA_64to4[4]                      = RX_DATA_6_net_2[4:4];
assign LANE_2_IOD_DQ_RX_DATA_65to5[5]                      = RX_DATA_6_net_2[5:5];
assign LANE_2_IOD_DQ_RX_DATA_66to6[6]                      = RX_DATA_6_net_2[6:6];
assign LANE_2_IOD_DQ_RX_DATA_67to7[7]                      = RX_DATA_6_net_2[7:7];
assign LANE_2_IOD_DQ_RX_DATA_70to0[0]                      = RX_DATA_7_net_2[0:0];
assign LANE_2_IOD_DQ_RX_DATA_71to1[1]                      = RX_DATA_7_net_2[1:1];
assign LANE_2_IOD_DQ_RX_DATA_72to2[2]                      = RX_DATA_7_net_2[2:2];
assign LANE_2_IOD_DQ_RX_DATA_73to3[3]                      = RX_DATA_7_net_2[3:3];
assign LANE_2_IOD_DQ_RX_DATA_74to4[4]                      = RX_DATA_7_net_2[4:4];
assign LANE_2_IOD_DQ_RX_DATA_75to5[5]                      = RX_DATA_7_net_2[5:5];
assign LANE_2_IOD_DQ_RX_DATA_76to6[6]                      = RX_DATA_7_net_2[6:6];
assign LANE_2_IOD_DQ_RX_DATA_77to7[7]                      = RX_DATA_7_net_2[7:7];
assign LANE_2_IOD_DQSW_TRAINING_RX_DATA_00to0[0]           = RX_DATA_0_net_10[0:0];
assign LANE_2_IOD_DQSW_TRAINING_RX_DATA_01to1[1]           = RX_DATA_0_net_10[1:1];
assign LANE_2_IOD_READ_TRAINING_RX_DATA_06to6[6]           = RX_DATA_0_net_11[6:6];
assign LANE_2_IOD_READ_TRAINING_RX_DATA_07to7[7]           = RX_DATA_0_net_11[7:7];
assign LANE_3_IOD_DQ_RX_DATA_00to0[0]                      = RX_DATA_0_net_12[0:0];
assign LANE_3_IOD_DQ_RX_DATA_01to1[1]                      = RX_DATA_0_net_12[1:1];
assign LANE_3_IOD_DQ_RX_DATA_02to2[2]                      = RX_DATA_0_net_12[2:2];
assign LANE_3_IOD_DQ_RX_DATA_03to3[3]                      = RX_DATA_0_net_12[3:3];
assign LANE_3_IOD_DQ_RX_DATA_04to4[4]                      = RX_DATA_0_net_12[4:4];
assign LANE_3_IOD_DQ_RX_DATA_05to5[5]                      = RX_DATA_0_net_12[5:5];
assign LANE_3_IOD_DQ_RX_DATA_06to6[6]                      = RX_DATA_0_net_12[6:6];
assign LANE_3_IOD_DQ_RX_DATA_07to7[7]                      = RX_DATA_0_net_12[7:7];
assign LANE_3_IOD_DQ_RX_DATA_10to0[0]                      = RX_DATA_1_net_3[0:0];
assign LANE_3_IOD_DQ_RX_DATA_11to1[1]                      = RX_DATA_1_net_3[1:1];
assign LANE_3_IOD_DQ_RX_DATA_12to2[2]                      = RX_DATA_1_net_3[2:2];
assign LANE_3_IOD_DQ_RX_DATA_13to3[3]                      = RX_DATA_1_net_3[3:3];
assign LANE_3_IOD_DQ_RX_DATA_14to4[4]                      = RX_DATA_1_net_3[4:4];
assign LANE_3_IOD_DQ_RX_DATA_15to5[5]                      = RX_DATA_1_net_3[5:5];
assign LANE_3_IOD_DQ_RX_DATA_16to6[6]                      = RX_DATA_1_net_3[6:6];
assign LANE_3_IOD_DQ_RX_DATA_17to7[7]                      = RX_DATA_1_net_3[7:7];
assign LANE_3_IOD_DQ_RX_DATA_20to0[0]                      = RX_DATA_2_net_3[0:0];
assign LANE_3_IOD_DQ_RX_DATA_21to1[1]                      = RX_DATA_2_net_3[1:1];
assign LANE_3_IOD_DQ_RX_DATA_22to2[2]                      = RX_DATA_2_net_3[2:2];
assign LANE_3_IOD_DQ_RX_DATA_23to3[3]                      = RX_DATA_2_net_3[3:3];
assign LANE_3_IOD_DQ_RX_DATA_24to4[4]                      = RX_DATA_2_net_3[4:4];
assign LANE_3_IOD_DQ_RX_DATA_25to5[5]                      = RX_DATA_2_net_3[5:5];
assign LANE_3_IOD_DQ_RX_DATA_26to6[6]                      = RX_DATA_2_net_3[6:6];
assign LANE_3_IOD_DQ_RX_DATA_27to7[7]                      = RX_DATA_2_net_3[7:7];
assign LANE_3_IOD_DQ_RX_DATA_30to0[0]                      = RX_DATA_3_net_3[0:0];
assign LANE_3_IOD_DQ_RX_DATA_31to1[1]                      = RX_DATA_3_net_3[1:1];
assign LANE_3_IOD_DQ_RX_DATA_32to2[2]                      = RX_DATA_3_net_3[2:2];
assign LANE_3_IOD_DQ_RX_DATA_33to3[3]                      = RX_DATA_3_net_3[3:3];
assign LANE_3_IOD_DQ_RX_DATA_34to4[4]                      = RX_DATA_3_net_3[4:4];
assign LANE_3_IOD_DQ_RX_DATA_35to5[5]                      = RX_DATA_3_net_3[5:5];
assign LANE_3_IOD_DQ_RX_DATA_36to6[6]                      = RX_DATA_3_net_3[6:6];
assign LANE_3_IOD_DQ_RX_DATA_37to7[7]                      = RX_DATA_3_net_3[7:7];
assign LANE_3_IOD_DQ_RX_DATA_40to0[0]                      = RX_DATA_4_net_3[0:0];
assign LANE_3_IOD_DQ_RX_DATA_41to1[1]                      = RX_DATA_4_net_3[1:1];
assign LANE_3_IOD_DQ_RX_DATA_42to2[2]                      = RX_DATA_4_net_3[2:2];
assign LANE_3_IOD_DQ_RX_DATA_43to3[3]                      = RX_DATA_4_net_3[3:3];
assign LANE_3_IOD_DQ_RX_DATA_44to4[4]                      = RX_DATA_4_net_3[4:4];
assign LANE_3_IOD_DQ_RX_DATA_45to5[5]                      = RX_DATA_4_net_3[5:5];
assign LANE_3_IOD_DQ_RX_DATA_46to6[6]                      = RX_DATA_4_net_3[6:6];
assign LANE_3_IOD_DQ_RX_DATA_47to7[7]                      = RX_DATA_4_net_3[7:7];
assign LANE_3_IOD_DQ_RX_DATA_50to0[0]                      = RX_DATA_5_net_3[0:0];
assign LANE_3_IOD_DQ_RX_DATA_51to1[1]                      = RX_DATA_5_net_3[1:1];
assign LANE_3_IOD_DQ_RX_DATA_52to2[2]                      = RX_DATA_5_net_3[2:2];
assign LANE_3_IOD_DQ_RX_DATA_53to3[3]                      = RX_DATA_5_net_3[3:3];
assign LANE_3_IOD_DQ_RX_DATA_54to4[4]                      = RX_DATA_5_net_3[4:4];
assign LANE_3_IOD_DQ_RX_DATA_55to5[5]                      = RX_DATA_5_net_3[5:5];
assign LANE_3_IOD_DQ_RX_DATA_56to6[6]                      = RX_DATA_5_net_3[6:6];
assign LANE_3_IOD_DQ_RX_DATA_57to7[7]                      = RX_DATA_5_net_3[7:7];
assign LANE_3_IOD_DQ_RX_DATA_60to0[0]                      = RX_DATA_6_net_3[0:0];
assign LANE_3_IOD_DQ_RX_DATA_61to1[1]                      = RX_DATA_6_net_3[1:1];
assign LANE_3_IOD_DQ_RX_DATA_62to2[2]                      = RX_DATA_6_net_3[2:2];
assign LANE_3_IOD_DQ_RX_DATA_63to3[3]                      = RX_DATA_6_net_3[3:3];
assign LANE_3_IOD_DQ_RX_DATA_64to4[4]                      = RX_DATA_6_net_3[4:4];
assign LANE_3_IOD_DQ_RX_DATA_65to5[5]                      = RX_DATA_6_net_3[5:5];
assign LANE_3_IOD_DQ_RX_DATA_66to6[6]                      = RX_DATA_6_net_3[6:6];
assign LANE_3_IOD_DQ_RX_DATA_67to7[7]                      = RX_DATA_6_net_3[7:7];
assign LANE_3_IOD_DQ_RX_DATA_70to0[0]                      = RX_DATA_7_net_3[0:0];
assign LANE_3_IOD_DQ_RX_DATA_71to1[1]                      = RX_DATA_7_net_3[1:1];
assign LANE_3_IOD_DQ_RX_DATA_72to2[2]                      = RX_DATA_7_net_3[2:2];
assign LANE_3_IOD_DQ_RX_DATA_73to3[3]                      = RX_DATA_7_net_3[3:3];
assign LANE_3_IOD_DQ_RX_DATA_74to4[4]                      = RX_DATA_7_net_3[4:4];
assign LANE_3_IOD_DQ_RX_DATA_75to5[5]                      = RX_DATA_7_net_3[5:5];
assign LANE_3_IOD_DQ_RX_DATA_76to6[6]                      = RX_DATA_7_net_3[6:6];
assign LANE_3_IOD_DQ_RX_DATA_77to7[7]                      = RX_DATA_7_net_3[7:7];
assign LANE_3_IOD_DQSW_TRAINING_RX_DATA_00to0[0]           = RX_DATA_0_net_13[0:0];
assign LANE_3_IOD_DQSW_TRAINING_RX_DATA_01to1[1]           = RX_DATA_0_net_13[1:1];
assign LANE_3_IOD_READ_TRAINING_RX_DATA_06to6[6]           = RX_DATA_0_net_14[6:6];
assign LANE_3_IOD_READ_TRAINING_RX_DATA_07to7[7]           = RX_DATA_0_net_14[7:7];
assign RX_DATA_0_slice_0[0]                                = RX_DATA_0_net_0[0:0];
assign RX_DATA_0_slice_1[1]                                = RX_DATA_0_net_0[1:1];
assign RX_DATA_0_slice_2[2]                                = RX_DATA_0_net_0[2:2];
assign RX_DATA_0_slice_3[1]                                = RX_DATA_0_net_1[1:1];
assign RX_DATA_0_slice_4[3]                                = RX_DATA_0_net_1[3:3];
assign RX_DATA_0_slice_5[5]                                = RX_DATA_0_net_1[5:5];
assign RX_DATA_0_slice_6[7]                                = RX_DATA_0_net_1[7:7];
assign RX_DATA_0_slice_7[0]                                = RX_DATA_0_net_2[0:0];
assign RX_DATA_0_slice_8[1]                                = RX_DATA_0_net_2[1:1];
assign RX_DATA_0_slice_9[2]                                = RX_DATA_0_net_2[2:2];
assign RX_DATA_0_slice_10[3]                               = RX_DATA_0_net_2[3:3];
assign RX_DATA_0_slice_11[4]                               = RX_DATA_0_net_2[4:4];
assign RX_DATA_0_slice_12[5]                               = RX_DATA_0_net_2[5:5];
assign RX_DATA_0_slice_13[7]                               = RX_DATA_0_net_2[7:7];
assign ODT_DYN_LANE_slice_0[0]                             = ODT_DYN_LANE_net_0[0:0];
assign ODT_DYN_LANE_slice_1[1]                             = ODT_DYN_LANE_net_0[1:1];
assign ODT_DYN_LANE_slice_2[2]                             = ODT_DYN_LANE_net_0[2:2];
assign ODT_DYN_LANE_slice_3[3]                             = ODT_DYN_LANE_net_0[3:3];
assign IOG_WRDATA_MASK_P0_slice_0[0]                       = IOG_WRDATA_MASK_P0_net_0[0:0];
assign IOG_WRDATA_MASK_P0_slice_1[1]                       = IOG_WRDATA_MASK_P0_net_0[1:1];
assign IOG_WRDATA_MASK_P0_slice_2[2]                       = IOG_WRDATA_MASK_P0_net_0[2:2];
assign IOG_WRDATA_MASK_P0_slice_3[3]                       = IOG_WRDATA_MASK_P0_net_0[3:3];
assign IOG_WRDATA_MASK_P0_slice_4[4]                       = IOG_WRDATA_MASK_P0_net_0[4:4];
assign IOG_WRDATA_MASK_P0_slice_5[5]                       = IOG_WRDATA_MASK_P0_net_0[5:5];
assign IOG_WRDATA_MASK_P0_slice_6[6]                       = IOG_WRDATA_MASK_P0_net_0[6:6];
assign IOG_WRDATA_MASK_P0_slice_7[7]                       = IOG_WRDATA_MASK_P0_net_0[7:7];
assign IOG_WRDATA_MASK_P1_slice_0[0]                       = IOG_WRDATA_MASK_P1_net_0[0:0];
assign IOG_WRDATA_MASK_P1_slice_1[1]                       = IOG_WRDATA_MASK_P1_net_0[1:1];
assign IOG_WRDATA_MASK_P1_slice_2[2]                       = IOG_WRDATA_MASK_P1_net_0[2:2];
assign IOG_WRDATA_MASK_P1_slice_3[3]                       = IOG_WRDATA_MASK_P1_net_0[3:3];
assign IOG_WRDATA_MASK_P1_slice_4[4]                       = IOG_WRDATA_MASK_P1_net_0[4:4];
assign IOG_WRDATA_MASK_P1_slice_5[5]                       = IOG_WRDATA_MASK_P1_net_0[5:5];
assign IOG_WRDATA_MASK_P1_slice_6[6]                       = IOG_WRDATA_MASK_P1_net_0[6:6];
assign IOG_WRDATA_MASK_P1_slice_7[7]                       = IOG_WRDATA_MASK_P1_net_0[7:7];
assign IOG_WRDATA_MASK_P2_slice_0[0]                       = IOG_WRDATA_MASK_P2_net_0[0:0];
assign IOG_WRDATA_MASK_P2_slice_1[1]                       = IOG_WRDATA_MASK_P2_net_0[1:1];
assign IOG_WRDATA_MASK_P2_slice_2[2]                       = IOG_WRDATA_MASK_P2_net_0[2:2];
assign IOG_WRDATA_MASK_P2_slice_3[3]                       = IOG_WRDATA_MASK_P2_net_0[3:3];
assign IOG_WRDATA_MASK_P2_slice_4[4]                       = IOG_WRDATA_MASK_P2_net_0[4:4];
assign IOG_WRDATA_MASK_P2_slice_5[5]                       = IOG_WRDATA_MASK_P2_net_0[5:5];
assign IOG_WRDATA_MASK_P2_slice_6[6]                       = IOG_WRDATA_MASK_P2_net_0[6:6];
assign IOG_WRDATA_MASK_P2_slice_7[7]                       = IOG_WRDATA_MASK_P2_net_0[7:7];
assign IOG_WRDATA_MASK_P3_slice_0[0]                       = IOG_WRDATA_MASK_P3_net_0[0:0];
assign IOG_WRDATA_MASK_P3_slice_1[1]                       = IOG_WRDATA_MASK_P3_net_0[1:1];
assign IOG_WRDATA_MASK_P3_slice_2[2]                       = IOG_WRDATA_MASK_P3_net_0[2:2];
assign IOG_WRDATA_MASK_P3_slice_3[3]                       = IOG_WRDATA_MASK_P3_net_0[3:3];
assign IOG_WRDATA_MASK_P3_slice_4[4]                       = IOG_WRDATA_MASK_P3_net_0[4:4];
assign IOG_WRDATA_MASK_P3_slice_5[5]                       = IOG_WRDATA_MASK_P3_net_0[5:5];
assign IOG_WRDATA_MASK_P3_slice_6[6]                       = IOG_WRDATA_MASK_P3_net_0[6:6];
assign IOG_WRDATA_MASK_P3_slice_7[7]                       = IOG_WRDATA_MASK_P3_net_0[7:7];
assign IOG_ADDRESS_P0_slice_0[14]                          = IOG_ADDRESS_P0_net_0[14:14];
assign IOG_ADDRESS_P0_slice_1[15]                          = IOG_ADDRESS_P0_net_0[15:15];
assign IOG_ADDRESS_P0_slice_2[16]                          = IOG_ADDRESS_P0_net_0[16:16];
assign IOG_ADDRESS_P0_slice_3[17]                          = IOG_ADDRESS_P0_net_0[17:17];
assign IOG_ADDRESS_P0_slice_4[18]                          = IOG_ADDRESS_P0_net_0[18:18];
assign IOG_ADDRESS_P0_slice_5[19]                          = IOG_ADDRESS_P0_net_0[19:19];
assign IOG_ADDRESS_P1_slice_0[14]                          = IOG_ADDRESS_P1_net_0[14:14];
assign IOG_ADDRESS_P1_slice_1[15]                          = IOG_ADDRESS_P1_net_0[15:15];
assign IOG_ADDRESS_P1_slice_2[16]                          = IOG_ADDRESS_P1_net_0[16:16];
assign IOG_ADDRESS_P1_slice_3[17]                          = IOG_ADDRESS_P1_net_0[17:17];
assign IOG_ADDRESS_P1_slice_4[18]                          = IOG_ADDRESS_P1_net_0[18:18];
assign IOG_ADDRESS_P1_slice_5[19]                          = IOG_ADDRESS_P1_net_0[19:19];
assign IOG_ADDRESS_P2_slice_0[14]                          = IOG_ADDRESS_P2_net_0[14:14];
assign IOG_ADDRESS_P2_slice_1[15]                          = IOG_ADDRESS_P2_net_0[15:15];
assign IOG_ADDRESS_P2_slice_2[16]                          = IOG_ADDRESS_P2_net_0[16:16];
assign IOG_ADDRESS_P2_slice_3[17]                          = IOG_ADDRESS_P2_net_0[17:17];
assign IOG_ADDRESS_P2_slice_4[18]                          = IOG_ADDRESS_P2_net_0[18:18];
assign IOG_ADDRESS_P2_slice_5[19]                          = IOG_ADDRESS_P2_net_0[19:19];
assign IOG_ADDRESS_P3_slice_0[14]                          = IOG_ADDRESS_P3_net_0[14:14];
assign IOG_ADDRESS_P3_slice_1[15]                          = IOG_ADDRESS_P3_net_0[15:15];
assign IOG_ADDRESS_P3_slice_2[16]                          = IOG_ADDRESS_P3_net_0[16:16];
assign IOG_ADDRESS_P3_slice_3[17]                          = IOG_ADDRESS_P3_net_0[17:17];
assign IOG_ADDRESS_P3_slice_4[18]                          = IOG_ADDRESS_P3_net_0[18:18];
assign IOG_ADDRESS_P3_slice_5[19]                          = IOG_ADDRESS_P3_net_0[19:19];
assign DFI_BANK_P0_OUT_slice_0[2]                          = DFI_BANK_P0_OUT_net_0[2:2];
assign DFI_BANK_P1_OUT_slice_0[2]                          = DFI_BANK_P1_OUT_net_0[2:2];
assign DFI_BANK_P2_OUT_slice_0[2]                          = DFI_BANK_P2_OUT_net_0[2:2];
assign DFI_BANK_P3_OUT_slice_0[2]                          = DFI_BANK_P3_OUT_net_0[2:2];
assign RX_DATA_0_slice_14[0]                               = RX_DATA_0_net_5[0:0];
assign RX_DATA_0_slice_15[1]                               = RX_DATA_0_net_5[1:1];
assign RX_DATA_0_slice_16[2]                               = RX_DATA_0_net_5[2:2];
assign RX_DATA_0_slice_17[3]                               = RX_DATA_0_net_5[3:3];
assign RX_DATA_0_slice_18[4]                               = RX_DATA_0_net_5[4:4];
assign RX_DATA_0_slice_19[5]                               = RX_DATA_0_net_5[5:5];
assign RX_DATA_0_slice_20[0]                               = RX_DATA_0_net_8[0:0];
assign RX_DATA_0_slice_21[1]                               = RX_DATA_0_net_8[1:1];
assign RX_DATA_0_slice_22[2]                               = RX_DATA_0_net_8[2:2];
assign RX_DATA_0_slice_23[3]                               = RX_DATA_0_net_8[3:3];
assign RX_DATA_0_slice_24[4]                               = RX_DATA_0_net_8[4:4];
assign RX_DATA_0_slice_25[5]                               = RX_DATA_0_net_8[5:5];
assign RX_DATA_0_slice_26[0]                               = RX_DATA_0_net_11[0:0];
assign RX_DATA_0_slice_27[1]                               = RX_DATA_0_net_11[1:1];
assign RX_DATA_0_slice_28[2]                               = RX_DATA_0_net_11[2:2];
assign RX_DATA_0_slice_29[3]                               = RX_DATA_0_net_11[3:3];
assign RX_DATA_0_slice_30[4]                               = RX_DATA_0_net_11[4:4];
assign RX_DATA_0_slice_31[5]                               = RX_DATA_0_net_11[5:5];
assign RX_DATA_0_slice_32[0]                               = RX_DATA_0_net_14[0:0];
assign RX_DATA_0_slice_33[1]                               = RX_DATA_0_net_14[1:1];
assign RX_DATA_0_slice_34[2]                               = RX_DATA_0_net_14[2:2];
assign RX_DATA_0_slice_35[3]                               = RX_DATA_0_net_14[3:3];
assign RX_DATA_0_slice_36[4]                               = RX_DATA_0_net_14[4:4];
assign RX_DATA_0_slice_37[5]                               = RX_DATA_0_net_14[5:5];
//--------------------------------------------------------------------
// Concatenation assignments
//--------------------------------------------------------------------
assign TX_DATA_0_net_0                 = { IOD_TRAINING_0_IOG_ADDRESS_P30to0[0] , IOD_TRAINING_0_IOG_ADDRESS_P20to0[0] , IOD_TRAINING_0_IOG_ADDRESS_P10to0[0] , IOD_TRAINING_0_IOG_ADDRESS_P00to0[0] };
assign TX_DATA_1_net_0                 = { IOD_TRAINING_0_IOG_ADDRESS_P31to1[1] , IOD_TRAINING_0_IOG_ADDRESS_P21to1[1] , IOD_TRAINING_0_IOG_ADDRESS_P11to1[1] , IOD_TRAINING_0_IOG_ADDRESS_P01to1[1] };
assign TX_DATA_2_net_0                 = { IOD_TRAINING_0_IOG_ADDRESS_P32to2[2] , IOD_TRAINING_0_IOG_ADDRESS_P22to2[2] , IOD_TRAINING_0_IOG_ADDRESS_P12to2[2] , IOD_TRAINING_0_IOG_ADDRESS_P02to2[2] };
assign TX_DATA_3_net_0                 = { IOD_TRAINING_0_IOG_ADDRESS_P33to3[3] , IOD_TRAINING_0_IOG_ADDRESS_P23to3[3] , IOD_TRAINING_0_IOG_ADDRESS_P13to3[3] , IOD_TRAINING_0_IOG_ADDRESS_P03to3[3] };
assign TX_DATA_4_net_0                 = { IOD_TRAINING_0_IOG_ADDRESS_P34to4[4] , IOD_TRAINING_0_IOG_ADDRESS_P24to4[4] , IOD_TRAINING_0_IOG_ADDRESS_P14to4[4] , IOD_TRAINING_0_IOG_ADDRESS_P04to4[4] };
assign TX_DATA_5_net_0                 = { IOD_TRAINING_0_IOG_ADDRESS_P35to5[5] , IOD_TRAINING_0_IOG_ADDRESS_P25to5[5] , IOD_TRAINING_0_IOG_ADDRESS_P15to5[5] , IOD_TRAINING_0_IOG_ADDRESS_P05to5[5] };
assign TX_DATA_6_net_0                 = { IOD_TRAINING_0_IOG_ADDRESS_P36to6[6] , IOD_TRAINING_0_IOG_ADDRESS_P26to6[6] , IOD_TRAINING_0_IOG_ADDRESS_P16to6[6] , IOD_TRAINING_0_IOG_ADDRESS_P06to6[6] };
assign TX_DATA_7_net_0                 = { IOD_TRAINING_0_IOG_ADDRESS_P37to7[7] , IOD_TRAINING_0_IOG_ADDRESS_P27to7[7] , IOD_TRAINING_0_IOG_ADDRESS_P17to7[7] , IOD_TRAINING_0_IOG_ADDRESS_P07to7[7] };
assign TX_DATA_8_net_0                 = { IOD_TRAINING_0_IOG_ADDRESS_P38to8[8] , IOD_TRAINING_0_IOG_ADDRESS_P28to8[8] , IOD_TRAINING_0_IOG_ADDRESS_P18to8[8] , IOD_TRAINING_0_IOG_ADDRESS_P08to8[8] };
assign TX_DATA_9_net_0                 = { IOD_TRAINING_0_IOG_ADDRESS_P39to9[9] , IOD_TRAINING_0_IOG_ADDRESS_P29to9[9] , IOD_TRAINING_0_IOG_ADDRESS_P19to9[9] , IOD_TRAINING_0_IOG_ADDRESS_P09to9[9] };
assign TX_DATA_10_net_0                = { IOD_TRAINING_0_IOG_ADDRESS_P310to10[10] , IOD_TRAINING_0_IOG_ADDRESS_P210to10[10] , IOD_TRAINING_0_IOG_ADDRESS_P110to10[10] , IOD_TRAINING_0_IOG_ADDRESS_P010to10[10] };
assign TX_DATA_11_net_0                = { IOD_TRAINING_0_IOG_ADDRESS_P311to11[11] , IOD_TRAINING_0_IOG_ADDRESS_P211to11[11] , IOD_TRAINING_0_IOG_ADDRESS_P111to11[11] , IOD_TRAINING_0_IOG_ADDRESS_P011to11[11] };
assign TX_DATA_0_net_1                 = { IOD_TRAINING_0_IOG_ADDRESS_P312to12[12] , IOD_TRAINING_0_IOG_ADDRESS_P212to12[12] , IOD_TRAINING_0_IOG_ADDRESS_P112to12[12] , IOD_TRAINING_0_IOG_ADDRESS_P012to12[12] };
assign OE_DATA_0_net_0                 = { IOD_TRAINING_0_CMD_OE , IOD_TRAINING_0_CMD_OE , IOD_TRAINING_0_CMD_OE , IOD_TRAINING_0_CMD_OE };
assign TX_DATA_0_net_2                 = { IOD_TRAINING_0_IOG_ADDRESS_P313to13[13] , IOD_TRAINING_0_IOG_ADDRESS_P213to13[13] , IOD_TRAINING_0_IOG_ADDRESS_P113to13[13] , IOD_TRAINING_0_IOG_ADDRESS_P013to13[13] };
assign TX_DATA_0_net_3                 = { IOD_TRAINING_0_DFI_ACT_N_P3_OUT , IOD_TRAINING_0_DFI_ACT_N_P2_OUT , IOD_TRAINING_0_DFI_ACT_N_P1_OUT , IOD_TRAINING_0_DFI_ACT_N_P0_OUT };
assign TX_DATA_0_net_4                 = { IOD_TRAINING_0_DFI_BANK_P3_OUT0to0[0] , IOD_TRAINING_0_DFI_BANK_P2_OUT0to0[0] , IOD_TRAINING_0_DFI_BANK_P1_OUT0to0[0] , IOD_TRAINING_0_DFI_BANK_P0_OUT0to0[0] };
assign TX_DATA_1_net_1                 = { IOD_TRAINING_0_DFI_BANK_P3_OUT1to1[1] , IOD_TRAINING_0_DFI_BANK_P2_OUT1to1[1] , IOD_TRAINING_0_DFI_BANK_P1_OUT1to1[1] , IOD_TRAINING_0_DFI_BANK_P0_OUT1to1[1] };
assign TX_DATA_0_net_5                 = { IOD_TRAINING_0_DFI_BG_P3_OUT0to0[0] , IOD_TRAINING_0_DFI_BG_P2_OUT0to0[0] , IOD_TRAINING_0_DFI_BG_P1_OUT0to0[0] , IOD_TRAINING_0_DFI_BG_P0_OUT0to0[0] };
assign TX_DATA_1_net_2                 = { IOD_TRAINING_0_DFI_BG_P3_OUT1to1[1] , IOD_TRAINING_0_DFI_BG_P2_OUT1to1[1] , IOD_TRAINING_0_DFI_BG_P1_OUT1to1[1] , IOD_TRAINING_0_DFI_BG_P0_OUT1to1[1] };
assign TX_DATA_0_net_6                 = { IOD_TRAINING_0_DFI_CAS_N_P3_OUT , IOD_TRAINING_0_DFI_CAS_N_P2_OUT , IOD_TRAINING_0_DFI_CAS_N_P1_OUT , IOD_TRAINING_0_DFI_CAS_N_P0_OUT };
assign TX_DATA_0_net_7                 = { IOD_TRAINING_0_DFI_CKE_P3_OUT , IOD_TRAINING_0_DFI_CKE_P2_OUT , IOD_TRAINING_0_DFI_CKE_P1_OUT , IOD_TRAINING_0_DFI_CKE_P0_OUT };
assign TX_DATA_0_net_8                 = { IOD_TRAINING_0_DFI_CS_N_P3_OUT , IOD_TRAINING_0_DFI_CS_N_P2_OUT , IOD_TRAINING_0_DFI_CS_N_P1_OUT , IOD_TRAINING_0_DFI_CS_N_P0_OUT };
assign TX_DATA_0_net_9                 = { IOD_TRAINING_0_DFI_ODT_P3_OUT , IOD_TRAINING_0_DFI_ODT_P2_OUT , IOD_TRAINING_0_DFI_ODT_P1_OUT , IOD_TRAINING_0_DFI_ODT_P0_OUT };
assign TX_DATA_0_net_10                = { IOD_TRAINING_0_DFI_RAS_N_P3_OUT , IOD_TRAINING_0_DFI_RAS_N_P2_OUT , IOD_TRAINING_0_DFI_RAS_N_P1_OUT , IOD_TRAINING_0_DFI_RAS_N_P0_OUT };
assign TX_DATA_0_net_11                = { IOD_TRAINING_0_DFI_RESET_N_P3_OUT , IOD_TRAINING_0_DFI_RESET_N_P2_OUT , IOD_TRAINING_0_DFI_RESET_N_P1_OUT , IOD_TRAINING_0_DFI_RESET_N_P0_OUT };
assign TX_DATA_0_net_12                = { IOD_TRAINING_0_DFI_WE_N_P3_OUT , IOD_TRAINING_0_DFI_WE_N_P2_OUT , IOD_TRAINING_0_DFI_WE_N_P1_OUT , IOD_TRAINING_0_DFI_WE_N_P0_OUT };
assign HS_IO_CLK_net_0                 = { HS_IO_CLK_270 , HS_IO_CLK };
assign READ_CLK_SEL_net_0              = { IOD_TRAINING_0_CLK_SEL2to2[2] , IOD_TRAINING_0_CLK_SEL1to1[1] , IOD_TRAINING_0_CLK_SEL0to0[0] };
assign TX_DATA_0_net_13                = { IOD_TRAINING_0_IOG_DM_TXDATA_OUT7to7[7] , IOD_TRAINING_0_IOG_DM_TXDATA_OUT6to6[6] , IOD_TRAINING_0_IOG_DM_TXDATA_OUT5to5[5] , IOD_TRAINING_0_IOG_DM_TXDATA_OUT4to4[4] , IOD_TRAINING_0_IOG_DM_TXDATA_OUT3to3[3] , IOD_TRAINING_0_IOG_DM_TXDATA_OUT2to2[2] , IOD_TRAINING_0_IOG_DM_TXDATA_OUT1to1[1] , IOD_TRAINING_0_IOG_DM_TXDATA_OUT0to0[0] };
assign OE_DATA_0_net_1                 = { IOD_TRAINING_0_DM_OE_P30to0[0] , IOD_TRAINING_0_DM_OE_P20to0[0] , IOD_TRAINING_0_DM_OE_P10to0[0] , IOD_TRAINING_0_DM_OE_P00to0[0] };
assign TX_DATA_0_net_14                = { IOD_TRAINING_0_IOG_DQ_TXDATA_OUT7to7[7] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT6to6[6] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT5to5[5] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT4to4[4] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT3to3[3] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT2to2[2] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT1to1[1] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT0to0[0] };
assign TX_DATA_1_net_3                 = { IOD_TRAINING_0_IOG_DQ_TXDATA_OUT15to15[15] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT14to14[14] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT13to13[13] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT12to12[12] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT11to11[11] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT10to10[10] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT9to9[9] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT8to8[8] };
assign TX_DATA_2_net_1                 = { IOD_TRAINING_0_IOG_DQ_TXDATA_OUT23to23[23] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT22to22[22] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT21to21[21] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT20to20[20] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT19to19[19] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT18to18[18] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT17to17[17] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT16to16[16] };
assign TX_DATA_3_net_1                 = { IOD_TRAINING_0_IOG_DQ_TXDATA_OUT31to31[31] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT30to30[30] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT29to29[29] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT28to28[28] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT27to27[27] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT26to26[26] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT25to25[25] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT24to24[24] };
assign TX_DATA_4_net_1                 = { IOD_TRAINING_0_IOG_DQ_TXDATA_OUT39to39[39] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT38to38[38] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT37to37[37] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT36to36[36] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT35to35[35] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT34to34[34] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT33to33[33] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT32to32[32] };
assign TX_DATA_5_net_1                 = { IOD_TRAINING_0_IOG_DQ_TXDATA_OUT47to47[47] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT46to46[46] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT45to45[45] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT44to44[44] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT43to43[43] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT42to42[42] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT41to41[41] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT40to40[40] };
assign TX_DATA_6_net_1                 = { IOD_TRAINING_0_IOG_DQ_TXDATA_OUT55to55[55] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT54to54[54] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT53to53[53] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT52to52[52] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT51to51[51] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT50to50[50] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT49to49[49] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT48to48[48] };
assign TX_DATA_7_net_1                 = { IOD_TRAINING_0_IOG_DQ_TXDATA_OUT63to63[63] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT62to62[62] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT61to61[61] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT60to60[60] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT59to59[59] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT58to58[58] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT57to57[57] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT56to56[56] };
assign OE_DATA_0_net_2                 = { IOD_TRAINING_0_IOG_OE_P30to0[0] , IOD_TRAINING_0_IOG_OE_P20to0[0] , IOD_TRAINING_0_IOG_OE_P10to0[0] , IOD_TRAINING_0_IOG_OE_P00to0[0] };
assign OE_DATA_1_net_0                 = { IOD_TRAINING_0_IOG_OE_P30to0[0] , IOD_TRAINING_0_IOG_OE_P20to0[0] , IOD_TRAINING_0_IOG_OE_P10to0[0] , IOD_TRAINING_0_IOG_OE_P00to0[0] };
assign OE_DATA_2_net_0                 = { IOD_TRAINING_0_IOG_OE_P30to0[0] , IOD_TRAINING_0_IOG_OE_P20to0[0] , IOD_TRAINING_0_IOG_OE_P10to0[0] , IOD_TRAINING_0_IOG_OE_P00to0[0] };
assign OE_DATA_3_net_0                 = { IOD_TRAINING_0_IOG_OE_P30to0[0] , IOD_TRAINING_0_IOG_OE_P20to0[0] , IOD_TRAINING_0_IOG_OE_P10to0[0] , IOD_TRAINING_0_IOG_OE_P00to0[0] };
assign OE_DATA_4_net_0                 = { IOD_TRAINING_0_IOG_OE_P30to0[0] , IOD_TRAINING_0_IOG_OE_P20to0[0] , IOD_TRAINING_0_IOG_OE_P10to0[0] , IOD_TRAINING_0_IOG_OE_P00to0[0] };
assign OE_DATA_5_net_0                 = { IOD_TRAINING_0_IOG_OE_P30to0[0] , IOD_TRAINING_0_IOG_OE_P20to0[0] , IOD_TRAINING_0_IOG_OE_P10to0[0] , IOD_TRAINING_0_IOG_OE_P00to0[0] };
assign OE_DATA_6_net_0                 = { IOD_TRAINING_0_IOG_OE_P30to0[0] , IOD_TRAINING_0_IOG_OE_P20to0[0] , IOD_TRAINING_0_IOG_OE_P10to0[0] , IOD_TRAINING_0_IOG_OE_P00to0[0] };
assign OE_DATA_7_net_0                 = { IOD_TRAINING_0_IOG_OE_P30to0[0] , IOD_TRAINING_0_IOG_OE_P20to0[0] , IOD_TRAINING_0_IOG_OE_P10to0[0] , IOD_TRAINING_0_IOG_OE_P00to0[0] };
assign OE_DATA_0_net_3                 = { IOD_TRAINING_0_DQS_OE_P30to0[0] , IOD_TRAINING_0_DQS_OE_P20to0[0] , IOD_TRAINING_0_DQS_OE_P10to0[0] , IOD_TRAINING_0_DQS_OE_P00to0[0] };
assign TX_DATA_0_net_15                = { IOD_TRAINING_0_IOG_RDDATA_EN_P3_N0to0[0] , IOD_TRAINING_0_IOG_RDDATA_EN_P3_P0to0[0] , IOD_TRAINING_0_IOG_RDDATA_EN_P2_N0to0[0] , IOD_TRAINING_0_IOG_RDDATA_EN_P2_P0to0[0] , IOD_TRAINING_0_IOG_RDDATA_EN_P1_N0to0[0] , IOD_TRAINING_0_IOG_RDDATA_EN_P1_P0to0[0] , IOD_TRAINING_0_IOG_RDDATA_EN_P0_N0to0[0] , IOD_TRAINING_0_IOG_RDDATA_EN_P0_P0to0[0] };
assign OE_DATA_0_net_4                 = { DFI_INIT_COMPLETE_net_0 , DFI_INIT_COMPLETE_net_0 , DFI_INIT_COMPLETE_net_0 , DFI_INIT_COMPLETE_net_0 };
assign HS_IO_CLK_net_1                 = { HS_IO_CLK_270 , HS_IO_CLK };
assign READ_CLK_SEL_net_1              = { IOD_TRAINING_0_CLK_SEL5to5[5] , IOD_TRAINING_0_CLK_SEL4to4[4] , IOD_TRAINING_0_CLK_SEL3to3[3] };
assign TX_DATA_0_net_16                = { IOD_TRAINING_0_IOG_DM_TXDATA_OUT15to15[15] , IOD_TRAINING_0_IOG_DM_TXDATA_OUT14to14[14] , IOD_TRAINING_0_IOG_DM_TXDATA_OUT13to13[13] , IOD_TRAINING_0_IOG_DM_TXDATA_OUT12to12[12] , IOD_TRAINING_0_IOG_DM_TXDATA_OUT11to11[11] , IOD_TRAINING_0_IOG_DM_TXDATA_OUT10to10[10] , IOD_TRAINING_0_IOG_DM_TXDATA_OUT9to9[9] , IOD_TRAINING_0_IOG_DM_TXDATA_OUT8to8[8] };
assign OE_DATA_0_net_5                 = { IOD_TRAINING_0_DM_OE_P31to1[1] , IOD_TRAINING_0_DM_OE_P21to1[1] , IOD_TRAINING_0_DM_OE_P11to1[1] , IOD_TRAINING_0_DM_OE_P01to1[1] };
assign TX_DATA_0_net_17                = { IOD_TRAINING_0_IOG_DQ_TXDATA_OUT71to71[71] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT70to70[70] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT69to69[69] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT68to68[68] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT67to67[67] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT66to66[66] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT65to65[65] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT64to64[64] };
assign TX_DATA_1_net_4                 = { IOD_TRAINING_0_IOG_DQ_TXDATA_OUT79to79[79] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT78to78[78] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT77to77[77] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT76to76[76] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT75to75[75] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT74to74[74] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT73to73[73] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT72to72[72] };
assign TX_DATA_2_net_2                 = { IOD_TRAINING_0_IOG_DQ_TXDATA_OUT87to87[87] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT86to86[86] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT85to85[85] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT84to84[84] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT83to83[83] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT82to82[82] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT81to81[81] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT80to80[80] };
assign TX_DATA_3_net_2                 = { IOD_TRAINING_0_IOG_DQ_TXDATA_OUT95to95[95] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT94to94[94] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT93to93[93] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT92to92[92] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT91to91[91] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT90to90[90] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT89to89[89] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT88to88[88] };
assign TX_DATA_4_net_2                 = { IOD_TRAINING_0_IOG_DQ_TXDATA_OUT103to103[103] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT102to102[102] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT101to101[101] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT100to100[100] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT99to99[99] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT98to98[98] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT97to97[97] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT96to96[96] };
assign TX_DATA_5_net_2                 = { IOD_TRAINING_0_IOG_DQ_TXDATA_OUT111to111[111] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT110to110[110] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT109to109[109] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT108to108[108] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT107to107[107] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT106to106[106] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT105to105[105] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT104to104[104] };
assign TX_DATA_6_net_2                 = { IOD_TRAINING_0_IOG_DQ_TXDATA_OUT119to119[119] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT118to118[118] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT117to117[117] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT116to116[116] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT115to115[115] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT114to114[114] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT113to113[113] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT112to112[112] };
assign TX_DATA_7_net_2                 = { IOD_TRAINING_0_IOG_DQ_TXDATA_OUT127to127[127] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT126to126[126] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT125to125[125] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT124to124[124] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT123to123[123] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT122to122[122] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT121to121[121] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT120to120[120] };
assign OE_DATA_0_net_6                 = { IOD_TRAINING_0_IOG_OE_P31to1[1] , IOD_TRAINING_0_IOG_OE_P21to1[1] , IOD_TRAINING_0_IOG_OE_P11to1[1] , IOD_TRAINING_0_IOG_OE_P01to1[1] };
assign OE_DATA_1_net_1                 = { IOD_TRAINING_0_IOG_OE_P31to1[1] , IOD_TRAINING_0_IOG_OE_P21to1[1] , IOD_TRAINING_0_IOG_OE_P11to1[1] , IOD_TRAINING_0_IOG_OE_P01to1[1] };
assign OE_DATA_2_net_1                 = { IOD_TRAINING_0_IOG_OE_P31to1[1] , IOD_TRAINING_0_IOG_OE_P21to1[1] , IOD_TRAINING_0_IOG_OE_P11to1[1] , IOD_TRAINING_0_IOG_OE_P01to1[1] };
assign OE_DATA_3_net_1                 = { IOD_TRAINING_0_IOG_OE_P31to1[1] , IOD_TRAINING_0_IOG_OE_P21to1[1] , IOD_TRAINING_0_IOG_OE_P11to1[1] , IOD_TRAINING_0_IOG_OE_P01to1[1] };
assign OE_DATA_4_net_1                 = { IOD_TRAINING_0_IOG_OE_P31to1[1] , IOD_TRAINING_0_IOG_OE_P21to1[1] , IOD_TRAINING_0_IOG_OE_P11to1[1] , IOD_TRAINING_0_IOG_OE_P01to1[1] };
assign OE_DATA_5_net_1                 = { IOD_TRAINING_0_IOG_OE_P31to1[1] , IOD_TRAINING_0_IOG_OE_P21to1[1] , IOD_TRAINING_0_IOG_OE_P11to1[1] , IOD_TRAINING_0_IOG_OE_P01to1[1] };
assign OE_DATA_6_net_1                 = { IOD_TRAINING_0_IOG_OE_P31to1[1] , IOD_TRAINING_0_IOG_OE_P21to1[1] , IOD_TRAINING_0_IOG_OE_P11to1[1] , IOD_TRAINING_0_IOG_OE_P01to1[1] };
assign OE_DATA_7_net_1                 = { IOD_TRAINING_0_IOG_OE_P31to1[1] , IOD_TRAINING_0_IOG_OE_P21to1[1] , IOD_TRAINING_0_IOG_OE_P11to1[1] , IOD_TRAINING_0_IOG_OE_P01to1[1] };
assign OE_DATA_0_net_7                 = { IOD_TRAINING_0_DQS_OE_P31to1[1] , IOD_TRAINING_0_DQS_OE_P21to1[1] , IOD_TRAINING_0_DQS_OE_P11to1[1] , IOD_TRAINING_0_DQS_OE_P01to1[1] };
assign TX_DATA_0_net_18                = { IOD_TRAINING_0_IOG_RDDATA_EN_P3_N1to1[1] , IOD_TRAINING_0_IOG_RDDATA_EN_P3_P1to1[1] , IOD_TRAINING_0_IOG_RDDATA_EN_P2_N1to1[1] , IOD_TRAINING_0_IOG_RDDATA_EN_P2_P1to1[1] , IOD_TRAINING_0_IOG_RDDATA_EN_P1_N1to1[1] , IOD_TRAINING_0_IOG_RDDATA_EN_P1_P1to1[1] , IOD_TRAINING_0_IOG_RDDATA_EN_P0_N1to1[1] , IOD_TRAINING_0_IOG_RDDATA_EN_P0_P1to1[1] };
assign OE_DATA_0_net_8                 = { DFI_INIT_COMPLETE_net_0 , DFI_INIT_COMPLETE_net_0 , DFI_INIT_COMPLETE_net_0 , DFI_INIT_COMPLETE_net_0 };
assign HS_IO_CLK_net_2                 = { HS_IO_CLK_270 , HS_IO_CLK };
assign READ_CLK_SEL_net_2              = { IOD_TRAINING_0_CLK_SEL8to8[8] , IOD_TRAINING_0_CLK_SEL7to7[7] , IOD_TRAINING_0_CLK_SEL6to6[6] };
assign TX_DATA_0_net_19                = { IOD_TRAINING_0_IOG_DM_TXDATA_OUT23to23[23] , IOD_TRAINING_0_IOG_DM_TXDATA_OUT22to22[22] , IOD_TRAINING_0_IOG_DM_TXDATA_OUT21to21[21] , IOD_TRAINING_0_IOG_DM_TXDATA_OUT20to20[20] , IOD_TRAINING_0_IOG_DM_TXDATA_OUT19to19[19] , IOD_TRAINING_0_IOG_DM_TXDATA_OUT18to18[18] , IOD_TRAINING_0_IOG_DM_TXDATA_OUT17to17[17] , IOD_TRAINING_0_IOG_DM_TXDATA_OUT16to16[16] };
assign OE_DATA_0_net_9                 = { IOD_TRAINING_0_DM_OE_P32to2[2] , IOD_TRAINING_0_DM_OE_P22to2[2] , IOD_TRAINING_0_DM_OE_P12to2[2] , IOD_TRAINING_0_DM_OE_P02to2[2] };
assign TX_DATA_0_net_20                = { IOD_TRAINING_0_IOG_DQ_TXDATA_OUT135to135[135] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT134to134[134] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT133to133[133] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT132to132[132] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT131to131[131] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT130to130[130] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT129to129[129] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT128to128[128] };
assign TX_DATA_1_net_5                 = { IOD_TRAINING_0_IOG_DQ_TXDATA_OUT143to143[143] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT142to142[142] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT141to141[141] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT140to140[140] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT139to139[139] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT138to138[138] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT137to137[137] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT136to136[136] };
assign TX_DATA_2_net_3                 = { IOD_TRAINING_0_IOG_DQ_TXDATA_OUT151to151[151] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT150to150[150] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT149to149[149] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT148to148[148] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT147to147[147] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT146to146[146] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT145to145[145] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT144to144[144] };
assign TX_DATA_3_net_3                 = { IOD_TRAINING_0_IOG_DQ_TXDATA_OUT159to159[159] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT158to158[158] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT157to157[157] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT156to156[156] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT155to155[155] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT154to154[154] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT153to153[153] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT152to152[152] };
assign TX_DATA_4_net_3                 = { IOD_TRAINING_0_IOG_DQ_TXDATA_OUT167to167[167] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT166to166[166] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT165to165[165] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT164to164[164] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT163to163[163] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT162to162[162] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT161to161[161] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT160to160[160] };
assign TX_DATA_5_net_3                 = { IOD_TRAINING_0_IOG_DQ_TXDATA_OUT175to175[175] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT174to174[174] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT173to173[173] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT172to172[172] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT171to171[171] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT170to170[170] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT169to169[169] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT168to168[168] };
assign TX_DATA_6_net_3                 = { IOD_TRAINING_0_IOG_DQ_TXDATA_OUT183to183[183] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT182to182[182] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT181to181[181] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT180to180[180] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT179to179[179] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT178to178[178] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT177to177[177] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT176to176[176] };
assign TX_DATA_7_net_3                 = { IOD_TRAINING_0_IOG_DQ_TXDATA_OUT191to191[191] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT190to190[190] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT189to189[189] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT188to188[188] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT187to187[187] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT186to186[186] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT185to185[185] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT184to184[184] };
assign OE_DATA_0_net_10                = { IOD_TRAINING_0_IOG_OE_P32to2[2] , IOD_TRAINING_0_IOG_OE_P22to2[2] , IOD_TRAINING_0_IOG_OE_P12to2[2] , IOD_TRAINING_0_IOG_OE_P02to2[2] };
assign OE_DATA_1_net_2                 = { IOD_TRAINING_0_IOG_OE_P32to2[2] , IOD_TRAINING_0_IOG_OE_P22to2[2] , IOD_TRAINING_0_IOG_OE_P12to2[2] , IOD_TRAINING_0_IOG_OE_P02to2[2] };
assign OE_DATA_2_net_2                 = { IOD_TRAINING_0_IOG_OE_P32to2[2] , IOD_TRAINING_0_IOG_OE_P22to2[2] , IOD_TRAINING_0_IOG_OE_P12to2[2] , IOD_TRAINING_0_IOG_OE_P02to2[2] };
assign OE_DATA_3_net_2                 = { IOD_TRAINING_0_IOG_OE_P32to2[2] , IOD_TRAINING_0_IOG_OE_P22to2[2] , IOD_TRAINING_0_IOG_OE_P12to2[2] , IOD_TRAINING_0_IOG_OE_P02to2[2] };
assign OE_DATA_4_net_2                 = { IOD_TRAINING_0_IOG_OE_P32to2[2] , IOD_TRAINING_0_IOG_OE_P22to2[2] , IOD_TRAINING_0_IOG_OE_P12to2[2] , IOD_TRAINING_0_IOG_OE_P02to2[2] };
assign OE_DATA_5_net_2                 = { IOD_TRAINING_0_IOG_OE_P32to2[2] , IOD_TRAINING_0_IOG_OE_P22to2[2] , IOD_TRAINING_0_IOG_OE_P12to2[2] , IOD_TRAINING_0_IOG_OE_P02to2[2] };
assign OE_DATA_6_net_2                 = { IOD_TRAINING_0_IOG_OE_P32to2[2] , IOD_TRAINING_0_IOG_OE_P22to2[2] , IOD_TRAINING_0_IOG_OE_P12to2[2] , IOD_TRAINING_0_IOG_OE_P02to2[2] };
assign OE_DATA_7_net_2                 = { IOD_TRAINING_0_IOG_OE_P32to2[2] , IOD_TRAINING_0_IOG_OE_P22to2[2] , IOD_TRAINING_0_IOG_OE_P12to2[2] , IOD_TRAINING_0_IOG_OE_P02to2[2] };
assign OE_DATA_0_net_11                = { IOD_TRAINING_0_DQS_OE_P32to2[2] , IOD_TRAINING_0_DQS_OE_P22to2[2] , IOD_TRAINING_0_DQS_OE_P12to2[2] , IOD_TRAINING_0_DQS_OE_P02to2[2] };
assign TX_DATA_0_net_21                = { IOD_TRAINING_0_IOG_RDDATA_EN_P3_N2to2[2] , IOD_TRAINING_0_IOG_RDDATA_EN_P3_P2to2[2] , IOD_TRAINING_0_IOG_RDDATA_EN_P2_N2to2[2] , IOD_TRAINING_0_IOG_RDDATA_EN_P2_P2to2[2] , IOD_TRAINING_0_IOG_RDDATA_EN_P1_N2to2[2] , IOD_TRAINING_0_IOG_RDDATA_EN_P1_P2to2[2] , IOD_TRAINING_0_IOG_RDDATA_EN_P0_N2to2[2] , IOD_TRAINING_0_IOG_RDDATA_EN_P0_P2to2[2] };
assign OE_DATA_0_net_12                = { DFI_INIT_COMPLETE_net_0 , DFI_INIT_COMPLETE_net_0 , DFI_INIT_COMPLETE_net_0 , DFI_INIT_COMPLETE_net_0 };
assign HS_IO_CLK_net_3                 = { HS_IO_CLK_270 , HS_IO_CLK };
assign READ_CLK_SEL_net_3              = { IOD_TRAINING_0_CLK_SEL11to11[11] , IOD_TRAINING_0_CLK_SEL10to10[10] , IOD_TRAINING_0_CLK_SEL9to9[9] };
assign TX_DATA_0_net_22                = { IOD_TRAINING_0_IOG_DM_TXDATA_OUT31to31[31] , IOD_TRAINING_0_IOG_DM_TXDATA_OUT30to30[30] , IOD_TRAINING_0_IOG_DM_TXDATA_OUT29to29[29] , IOD_TRAINING_0_IOG_DM_TXDATA_OUT28to28[28] , IOD_TRAINING_0_IOG_DM_TXDATA_OUT27to27[27] , IOD_TRAINING_0_IOG_DM_TXDATA_OUT26to26[26] , IOD_TRAINING_0_IOG_DM_TXDATA_OUT25to25[25] , IOD_TRAINING_0_IOG_DM_TXDATA_OUT24to24[24] };
assign OE_DATA_0_net_13                = { IOD_TRAINING_0_DM_OE_P33to3[3] , IOD_TRAINING_0_DM_OE_P23to3[3] , IOD_TRAINING_0_DM_OE_P13to3[3] , IOD_TRAINING_0_DM_OE_P03to3[3] };
assign TX_DATA_0_net_23                = { IOD_TRAINING_0_IOG_DQ_TXDATA_OUT199to199[199] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT198to198[198] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT197to197[197] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT196to196[196] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT195to195[195] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT194to194[194] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT193to193[193] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT192to192[192] };
assign TX_DATA_1_net_6                 = { IOD_TRAINING_0_IOG_DQ_TXDATA_OUT207to207[207] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT206to206[206] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT205to205[205] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT204to204[204] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT203to203[203] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT202to202[202] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT201to201[201] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT200to200[200] };
assign TX_DATA_2_net_4                 = { IOD_TRAINING_0_IOG_DQ_TXDATA_OUT215to215[215] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT214to214[214] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT213to213[213] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT212to212[212] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT211to211[211] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT210to210[210] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT209to209[209] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT208to208[208] };
assign TX_DATA_3_net_4                 = { IOD_TRAINING_0_IOG_DQ_TXDATA_OUT223to223[223] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT222to222[222] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT221to221[221] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT220to220[220] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT219to219[219] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT218to218[218] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT217to217[217] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT216to216[216] };
assign TX_DATA_4_net_4                 = { IOD_TRAINING_0_IOG_DQ_TXDATA_OUT231to231[231] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT230to230[230] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT229to229[229] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT228to228[228] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT227to227[227] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT226to226[226] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT225to225[225] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT224to224[224] };
assign TX_DATA_5_net_4                 = { IOD_TRAINING_0_IOG_DQ_TXDATA_OUT239to239[239] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT238to238[238] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT237to237[237] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT236to236[236] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT235to235[235] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT234to234[234] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT233to233[233] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT232to232[232] };
assign TX_DATA_6_net_4                 = { IOD_TRAINING_0_IOG_DQ_TXDATA_OUT247to247[247] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT246to246[246] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT245to245[245] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT244to244[244] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT243to243[243] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT242to242[242] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT241to241[241] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT240to240[240] };
assign TX_DATA_7_net_4                 = { IOD_TRAINING_0_IOG_DQ_TXDATA_OUT255to255[255] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT254to254[254] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT253to253[253] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT252to252[252] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT251to251[251] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT250to250[250] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT249to249[249] , IOD_TRAINING_0_IOG_DQ_TXDATA_OUT248to248[248] };
assign OE_DATA_0_net_14                = { IOD_TRAINING_0_IOG_OE_P33to3[3] , IOD_TRAINING_0_IOG_OE_P23to3[3] , IOD_TRAINING_0_IOG_OE_P13to3[3] , IOD_TRAINING_0_IOG_OE_P03to3[3] };
assign OE_DATA_1_net_3                 = { IOD_TRAINING_0_IOG_OE_P33to3[3] , IOD_TRAINING_0_IOG_OE_P23to3[3] , IOD_TRAINING_0_IOG_OE_P13to3[3] , IOD_TRAINING_0_IOG_OE_P03to3[3] };
assign OE_DATA_2_net_3                 = { IOD_TRAINING_0_IOG_OE_P33to3[3] , IOD_TRAINING_0_IOG_OE_P23to3[3] , IOD_TRAINING_0_IOG_OE_P13to3[3] , IOD_TRAINING_0_IOG_OE_P03to3[3] };
assign OE_DATA_3_net_3                 = { IOD_TRAINING_0_IOG_OE_P33to3[3] , IOD_TRAINING_0_IOG_OE_P23to3[3] , IOD_TRAINING_0_IOG_OE_P13to3[3] , IOD_TRAINING_0_IOG_OE_P03to3[3] };
assign OE_DATA_4_net_3                 = { IOD_TRAINING_0_IOG_OE_P33to3[3] , IOD_TRAINING_0_IOG_OE_P23to3[3] , IOD_TRAINING_0_IOG_OE_P13to3[3] , IOD_TRAINING_0_IOG_OE_P03to3[3] };
assign OE_DATA_5_net_3                 = { IOD_TRAINING_0_IOG_OE_P33to3[3] , IOD_TRAINING_0_IOG_OE_P23to3[3] , IOD_TRAINING_0_IOG_OE_P13to3[3] , IOD_TRAINING_0_IOG_OE_P03to3[3] };
assign OE_DATA_6_net_3                 = { IOD_TRAINING_0_IOG_OE_P33to3[3] , IOD_TRAINING_0_IOG_OE_P23to3[3] , IOD_TRAINING_0_IOG_OE_P13to3[3] , IOD_TRAINING_0_IOG_OE_P03to3[3] };
assign OE_DATA_7_net_3                 = { IOD_TRAINING_0_IOG_OE_P33to3[3] , IOD_TRAINING_0_IOG_OE_P23to3[3] , IOD_TRAINING_0_IOG_OE_P13to3[3] , IOD_TRAINING_0_IOG_OE_P03to3[3] };
assign OE_DATA_0_net_15                = { IOD_TRAINING_0_DQS_OE_P33to3[3] , IOD_TRAINING_0_DQS_OE_P23to3[3] , IOD_TRAINING_0_DQS_OE_P13to3[3] , IOD_TRAINING_0_DQS_OE_P03to3[3] };
assign TX_DATA_0_net_24                = { IOD_TRAINING_0_IOG_RDDATA_EN_P3_N3to3[3] , IOD_TRAINING_0_IOG_RDDATA_EN_P3_P3to3[3] , IOD_TRAINING_0_IOG_RDDATA_EN_P2_N3to3[3] , IOD_TRAINING_0_IOG_RDDATA_EN_P2_P3to3[3] , IOD_TRAINING_0_IOG_RDDATA_EN_P1_N3to3[3] , IOD_TRAINING_0_IOG_RDDATA_EN_P1_P3to3[3] , IOD_TRAINING_0_IOG_RDDATA_EN_P0_N3to3[3] , IOD_TRAINING_0_IOG_RDDATA_EN_P0_P3to3[3] };
assign OE_DATA_0_net_16                = { DFI_INIT_COMPLETE_net_0 , DFI_INIT_COMPLETE_net_0 , DFI_INIT_COMPLETE_net_0 , DFI_INIT_COMPLETE_net_0 };
assign BURST_DETECT_net_0              = { LANE_3_CTRL_RX_BURST_DETECT , LANE_2_CTRL_RX_BURST_DETECT , LANE_1_CTRL_RX_BURST_DETECT , LANE_0_CTRL_RX_BURST_DETECT };
assign RX_OUT_OF_RANGE_net_0           = { LANE_3_CTRL_RX_DELAY_LINE_OUT_OF_RANGE , LANE_3_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_7 , LANE_3_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_6 , LANE_3_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_5 , LANE_3_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_4 , LANE_3_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_3 , LANE_3_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_2 , LANE_3_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_1 , LANE_3_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_0 , LANE_2_CTRL_RX_DELAY_LINE_OUT_OF_RANGE , LANE_2_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_7 , LANE_2_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_6 , LANE_2_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_5 , LANE_2_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_4 , LANE_2_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_3 , LANE_2_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_2 , LANE_2_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_1 , LANE_2_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_0 , LANE_1_CTRL_RX_DELAY_LINE_OUT_OF_RANGE , LANE_1_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_7 , LANE_1_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_6 , LANE_1_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_5 , LANE_1_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_4 , LANE_1_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_3 , LANE_1_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_2 , LANE_1_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_1 , LANE_1_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_0 , LANE_0_CTRL_RX_DELAY_LINE_OUT_OF_RANGE , LANE_0_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_7 , LANE_0_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_6 , LANE_0_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_5 , LANE_0_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_4 , LANE_0_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_3 , LANE_0_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_2 , LANE_0_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_1 , LANE_0_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_0 };
assign TX_OUT_OF_RANGE_net_0           = { LANE_3_CTRL_TX_DELAY_LINE_OUT_OF_RANGE , LANE_3_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_7 , LANE_3_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_6 , LANE_3_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_5 , LANE_3_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_4 , LANE_3_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_3 , LANE_3_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_2 , LANE_3_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_1 , LANE_3_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_0 , LANE_2_CTRL_TX_DELAY_LINE_OUT_OF_RANGE , LANE_2_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_7 , LANE_2_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_6 , LANE_2_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_5 , LANE_2_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_4 , LANE_2_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_3 , LANE_2_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_2 , LANE_2_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_1 , LANE_2_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_0 , LANE_1_CTRL_TX_DELAY_LINE_OUT_OF_RANGE , LANE_1_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_7 , LANE_1_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_6 , LANE_1_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_5 , LANE_1_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_4 , LANE_1_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_3 , LANE_1_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_2 , LANE_1_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_1 , LANE_1_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_0 , LANE_0_CTRL_TX_DELAY_LINE_OUT_OF_RANGE , LANE_0_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_7 , LANE_0_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_6 , LANE_0_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_5 , LANE_0_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_4 , LANE_0_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_3 , LANE_0_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_2 , LANE_0_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_1 , LANE_0_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_0 };
assign IOG_RDDATA_net_0                = { LANE_3_IOD_DQ_RX_DATA_77to7[7] , LANE_3_IOD_DQ_RX_DATA_67to7[7] , LANE_3_IOD_DQ_RX_DATA_57to7[7] , LANE_3_IOD_DQ_RX_DATA_47to7[7] , LANE_3_IOD_DQ_RX_DATA_37to7[7] , LANE_3_IOD_DQ_RX_DATA_27to7[7] , LANE_3_IOD_DQ_RX_DATA_17to7[7] , LANE_3_IOD_DQ_RX_DATA_07to7[7] , LANE_2_IOD_DQ_RX_DATA_77to7[7] , LANE_2_IOD_DQ_RX_DATA_67to7[7] , LANE_2_IOD_DQ_RX_DATA_57to7[7] , LANE_2_IOD_DQ_RX_DATA_47to7[7] , LANE_2_IOD_DQ_RX_DATA_37to7[7] , LANE_2_IOD_DQ_RX_DATA_27to7[7] , LANE_2_IOD_DQ_RX_DATA_17to7[7] , LANE_2_IOD_DQ_RX_DATA_07to7[7] , LANE_1_IOD_DQ_RX_DATA_77to7[7] , LANE_1_IOD_DQ_RX_DATA_67to7[7] , LANE_1_IOD_DQ_RX_DATA_57to7[7] , LANE_1_IOD_DQ_RX_DATA_47to7[7] , LANE_1_IOD_DQ_RX_DATA_37to7[7] , LANE_1_IOD_DQ_RX_DATA_27to7[7] , LANE_1_IOD_DQ_RX_DATA_17to7[7] , LANE_1_IOD_DQ_RX_DATA_07to7[7] , LANE_0_IOD_DQ_RX_DATA_77to7[7] , LANE_0_IOD_DQ_RX_DATA_67to7[7] , LANE_0_IOD_DQ_RX_DATA_57to7[7] , LANE_0_IOD_DQ_RX_DATA_47to7[7] , LANE_0_IOD_DQ_RX_DATA_37to7[7] , LANE_0_IOD_DQ_RX_DATA_27to7[7] , LANE_0_IOD_DQ_RX_DATA_17to7[7] , LANE_0_IOD_DQ_RX_DATA_07to7[7] , LANE_3_IOD_DQ_RX_DATA_76to6[6] , LANE_3_IOD_DQ_RX_DATA_66to6[6] , LANE_3_IOD_DQ_RX_DATA_56to6[6] , LANE_3_IOD_DQ_RX_DATA_46to6[6] , LANE_3_IOD_DQ_RX_DATA_36to6[6] , LANE_3_IOD_DQ_RX_DATA_26to6[6] , LANE_3_IOD_DQ_RX_DATA_16to6[6] , LANE_3_IOD_DQ_RX_DATA_06to6[6] , LANE_2_IOD_DQ_RX_DATA_76to6[6] , LANE_2_IOD_DQ_RX_DATA_66to6[6] , LANE_2_IOD_DQ_RX_DATA_56to6[6] , LANE_2_IOD_DQ_RX_DATA_46to6[6] , LANE_2_IOD_DQ_RX_DATA_36to6[6] , LANE_2_IOD_DQ_RX_DATA_26to6[6] , LANE_2_IOD_DQ_RX_DATA_16to6[6] , LANE_2_IOD_DQ_RX_DATA_06to6[6] , LANE_1_IOD_DQ_RX_DATA_76to6[6] , LANE_1_IOD_DQ_RX_DATA_66to6[6] , LANE_1_IOD_DQ_RX_DATA_56to6[6] , LANE_1_IOD_DQ_RX_DATA_46to6[6] , LANE_1_IOD_DQ_RX_DATA_36to6[6] , LANE_1_IOD_DQ_RX_DATA_26to6[6] , LANE_1_IOD_DQ_RX_DATA_16to6[6] , LANE_1_IOD_DQ_RX_DATA_06to6[6] , LANE_0_IOD_DQ_RX_DATA_76to6[6] , LANE_0_IOD_DQ_RX_DATA_66to6[6] , LANE_0_IOD_DQ_RX_DATA_56to6[6] , LANE_0_IOD_DQ_RX_DATA_46to6[6] , LANE_0_IOD_DQ_RX_DATA_36to6[6] , LANE_0_IOD_DQ_RX_DATA_26to6[6] , LANE_0_IOD_DQ_RX_DATA_16to6[6] , LANE_0_IOD_DQ_RX_DATA_06to6[6] , LANE_3_IOD_DQ_RX_DATA_75to5[5] , LANE_3_IOD_DQ_RX_DATA_65to5[5] , LANE_3_IOD_DQ_RX_DATA_55to5[5] , LANE_3_IOD_DQ_RX_DATA_45to5[5] , LANE_3_IOD_DQ_RX_DATA_35to5[5] , LANE_3_IOD_DQ_RX_DATA_25to5[5] , LANE_3_IOD_DQ_RX_DATA_15to5[5] , LANE_3_IOD_DQ_RX_DATA_05to5[5] , LANE_2_IOD_DQ_RX_DATA_75to5[5] , LANE_2_IOD_DQ_RX_DATA_65to5[5] , LANE_2_IOD_DQ_RX_DATA_55to5[5] , LANE_2_IOD_DQ_RX_DATA_45to5[5] , LANE_2_IOD_DQ_RX_DATA_35to5[5] , LANE_2_IOD_DQ_RX_DATA_25to5[5] , LANE_2_IOD_DQ_RX_DATA_15to5[5] , LANE_2_IOD_DQ_RX_DATA_05to5[5] , LANE_1_IOD_DQ_RX_DATA_75to5[5] , LANE_1_IOD_DQ_RX_DATA_65to5[5] , LANE_1_IOD_DQ_RX_DATA_55to5[5] , LANE_1_IOD_DQ_RX_DATA_45to5[5] , LANE_1_IOD_DQ_RX_DATA_35to5[5] , LANE_1_IOD_DQ_RX_DATA_25to5[5] , LANE_1_IOD_DQ_RX_DATA_15to5[5] , LANE_1_IOD_DQ_RX_DATA_05to5[5] , LANE_0_IOD_DQ_RX_DATA_75to5[5] , LANE_0_IOD_DQ_RX_DATA_65to5[5] , LANE_0_IOD_DQ_RX_DATA_55to5[5] , LANE_0_IOD_DQ_RX_DATA_45to5[5] , LANE_0_IOD_DQ_RX_DATA_35to5[5] , LANE_0_IOD_DQ_RX_DATA_25to5[5] , LANE_0_IOD_DQ_RX_DATA_15to5[5] , LANE_0_IOD_DQ_RX_DATA_05to5[5] , LANE_3_IOD_DQ_RX_DATA_74to4[4] , LANE_3_IOD_DQ_RX_DATA_64to4[4] , LANE_3_IOD_DQ_RX_DATA_54to4[4] , LANE_3_IOD_DQ_RX_DATA_44to4[4] , LANE_3_IOD_DQ_RX_DATA_34to4[4] , LANE_3_IOD_DQ_RX_DATA_24to4[4] , LANE_3_IOD_DQ_RX_DATA_14to4[4] , LANE_3_IOD_DQ_RX_DATA_04to4[4] , LANE_2_IOD_DQ_RX_DATA_74to4[4] , LANE_2_IOD_DQ_RX_DATA_64to4[4] , LANE_2_IOD_DQ_RX_DATA_54to4[4] , LANE_2_IOD_DQ_RX_DATA_44to4[4] , LANE_2_IOD_DQ_RX_DATA_34to4[4] , LANE_2_IOD_DQ_RX_DATA_24to4[4] , LANE_2_IOD_DQ_RX_DATA_14to4[4] , LANE_2_IOD_DQ_RX_DATA_04to4[4] , LANE_1_IOD_DQ_RX_DATA_74to4[4] , LANE_1_IOD_DQ_RX_DATA_64to4[4] , LANE_1_IOD_DQ_RX_DATA_54to4[4] , LANE_1_IOD_DQ_RX_DATA_44to4[4] , LANE_1_IOD_DQ_RX_DATA_34to4[4] , LANE_1_IOD_DQ_RX_DATA_24to4[4] , LANE_1_IOD_DQ_RX_DATA_14to4[4] , LANE_1_IOD_DQ_RX_DATA_04to4[4] , LANE_0_IOD_DQ_RX_DATA_74to4[4] , LANE_0_IOD_DQ_RX_DATA_64to4[4] , LANE_0_IOD_DQ_RX_DATA_54to4[4] , LANE_0_IOD_DQ_RX_DATA_44to4[4] , LANE_0_IOD_DQ_RX_DATA_34to4[4] , LANE_0_IOD_DQ_RX_DATA_24to4[4] , LANE_0_IOD_DQ_RX_DATA_14to4[4] , LANE_0_IOD_DQ_RX_DATA_04to4[4] , LANE_3_IOD_DQ_RX_DATA_73to3[3] , LANE_3_IOD_DQ_RX_DATA_63to3[3] , LANE_3_IOD_DQ_RX_DATA_53to3[3] , LANE_3_IOD_DQ_RX_DATA_43to3[3] , LANE_3_IOD_DQ_RX_DATA_33to3[3] , LANE_3_IOD_DQ_RX_DATA_23to3[3] , LANE_3_IOD_DQ_RX_DATA_13to3[3] , LANE_3_IOD_DQ_RX_DATA_03to3[3] , LANE_2_IOD_DQ_RX_DATA_73to3[3] , LANE_2_IOD_DQ_RX_DATA_63to3[3] , LANE_2_IOD_DQ_RX_DATA_53to3[3] , LANE_2_IOD_DQ_RX_DATA_43to3[3] , LANE_2_IOD_DQ_RX_DATA_33to3[3] , LANE_2_IOD_DQ_RX_DATA_23to3[3] , LANE_2_IOD_DQ_RX_DATA_13to3[3] , LANE_2_IOD_DQ_RX_DATA_03to3[3] , LANE_1_IOD_DQ_RX_DATA_73to3[3] , LANE_1_IOD_DQ_RX_DATA_63to3[3] , LANE_1_IOD_DQ_RX_DATA_53to3[3] , LANE_1_IOD_DQ_RX_DATA_43to3[3] , LANE_1_IOD_DQ_RX_DATA_33to3[3] , LANE_1_IOD_DQ_RX_DATA_23to3[3] , LANE_1_IOD_DQ_RX_DATA_13to3[3] , LANE_1_IOD_DQ_RX_DATA_03to3[3] , LANE_0_IOD_DQ_RX_DATA_73to3[3] , LANE_0_IOD_DQ_RX_DATA_63to3[3] , LANE_0_IOD_DQ_RX_DATA_53to3[3] , LANE_0_IOD_DQ_RX_DATA_43to3[3] , LANE_0_IOD_DQ_RX_DATA_33to3[3] , LANE_0_IOD_DQ_RX_DATA_23to3[3] , LANE_0_IOD_DQ_RX_DATA_13to3[3] , LANE_0_IOD_DQ_RX_DATA_03to3[3] , LANE_3_IOD_DQ_RX_DATA_72to2[2] , LANE_3_IOD_DQ_RX_DATA_62to2[2] , LANE_3_IOD_DQ_RX_DATA_52to2[2] , LANE_3_IOD_DQ_RX_DATA_42to2[2] , LANE_3_IOD_DQ_RX_DATA_32to2[2] , LANE_3_IOD_DQ_RX_DATA_22to2[2] , LANE_3_IOD_DQ_RX_DATA_12to2[2] , LANE_3_IOD_DQ_RX_DATA_02to2[2] , LANE_2_IOD_DQ_RX_DATA_72to2[2] , LANE_2_IOD_DQ_RX_DATA_62to2[2] , LANE_2_IOD_DQ_RX_DATA_52to2[2] , LANE_2_IOD_DQ_RX_DATA_42to2[2] , LANE_2_IOD_DQ_RX_DATA_32to2[2] , LANE_2_IOD_DQ_RX_DATA_22to2[2] , LANE_2_IOD_DQ_RX_DATA_12to2[2] , LANE_2_IOD_DQ_RX_DATA_02to2[2] , LANE_1_IOD_DQ_RX_DATA_72to2[2] , LANE_1_IOD_DQ_RX_DATA_62to2[2] , LANE_1_IOD_DQ_RX_DATA_52to2[2] , LANE_1_IOD_DQ_RX_DATA_42to2[2] , LANE_1_IOD_DQ_RX_DATA_32to2[2] , LANE_1_IOD_DQ_RX_DATA_22to2[2] , LANE_1_IOD_DQ_RX_DATA_12to2[2] , LANE_1_IOD_DQ_RX_DATA_02to2[2] , LANE_0_IOD_DQ_RX_DATA_72to2[2] , LANE_0_IOD_DQ_RX_DATA_62to2[2] , LANE_0_IOD_DQ_RX_DATA_52to2[2] , LANE_0_IOD_DQ_RX_DATA_42to2[2] , LANE_0_IOD_DQ_RX_DATA_32to2[2] , LANE_0_IOD_DQ_RX_DATA_22to2[2] , LANE_0_IOD_DQ_RX_DATA_12to2[2] , LANE_0_IOD_DQ_RX_DATA_02to2[2] , LANE_3_IOD_DQ_RX_DATA_71to1[1] , LANE_3_IOD_DQ_RX_DATA_61to1[1] , LANE_3_IOD_DQ_RX_DATA_51to1[1] , LANE_3_IOD_DQ_RX_DATA_41to1[1] , LANE_3_IOD_DQ_RX_DATA_31to1[1] , LANE_3_IOD_DQ_RX_DATA_21to1[1] , LANE_3_IOD_DQ_RX_DATA_11to1[1] , LANE_3_IOD_DQ_RX_DATA_01to1[1] , LANE_2_IOD_DQ_RX_DATA_71to1[1] , LANE_2_IOD_DQ_RX_DATA_61to1[1] , LANE_2_IOD_DQ_RX_DATA_51to1[1] , LANE_2_IOD_DQ_RX_DATA_41to1[1] , LANE_2_IOD_DQ_RX_DATA_31to1[1] , LANE_2_IOD_DQ_RX_DATA_21to1[1] , LANE_2_IOD_DQ_RX_DATA_11to1[1] , LANE_2_IOD_DQ_RX_DATA_01to1[1] , LANE_1_IOD_DQ_RX_DATA_71to1[1] , LANE_1_IOD_DQ_RX_DATA_61to1[1] , LANE_1_IOD_DQ_RX_DATA_51to1[1] , LANE_1_IOD_DQ_RX_DATA_41to1[1] , LANE_1_IOD_DQ_RX_DATA_31to1[1] , LANE_1_IOD_DQ_RX_DATA_21to1[1] , LANE_1_IOD_DQ_RX_DATA_11to1[1] , LANE_1_IOD_DQ_RX_DATA_01to1[1] , LANE_0_IOD_DQ_RX_DATA_71to1[1] , LANE_0_IOD_DQ_RX_DATA_61to1[1] , LANE_0_IOD_DQ_RX_DATA_51to1[1] , LANE_0_IOD_DQ_RX_DATA_41to1[1] , LANE_0_IOD_DQ_RX_DATA_31to1[1] , LANE_0_IOD_DQ_RX_DATA_21to1[1] , LANE_0_IOD_DQ_RX_DATA_11to1[1] , LANE_0_IOD_DQ_RX_DATA_01to1[1] , LANE_3_IOD_DQ_RX_DATA_70to0[0] , LANE_3_IOD_DQ_RX_DATA_60to0[0] , LANE_3_IOD_DQ_RX_DATA_50to0[0] , LANE_3_IOD_DQ_RX_DATA_40to0[0] , LANE_3_IOD_DQ_RX_DATA_30to0[0] , LANE_3_IOD_DQ_RX_DATA_20to0[0] , LANE_3_IOD_DQ_RX_DATA_10to0[0] , LANE_3_IOD_DQ_RX_DATA_00to0[0] , LANE_2_IOD_DQ_RX_DATA_70to0[0] , LANE_2_IOD_DQ_RX_DATA_60to0[0] , LANE_2_IOD_DQ_RX_DATA_50to0[0] , LANE_2_IOD_DQ_RX_DATA_40to0[0] , LANE_2_IOD_DQ_RX_DATA_30to0[0] , LANE_2_IOD_DQ_RX_DATA_20to0[0] , LANE_2_IOD_DQ_RX_DATA_10to0[0] , LANE_2_IOD_DQ_RX_DATA_00to0[0] , LANE_1_IOD_DQ_RX_DATA_70to0[0] , LANE_1_IOD_DQ_RX_DATA_60to0[0] , LANE_1_IOD_DQ_RX_DATA_50to0[0] , LANE_1_IOD_DQ_RX_DATA_40to0[0] , LANE_1_IOD_DQ_RX_DATA_30to0[0] , LANE_1_IOD_DQ_RX_DATA_20to0[0] , LANE_1_IOD_DQ_RX_DATA_10to0[0] , LANE_1_IOD_DQ_RX_DATA_00to0[0] , LANE_0_IOD_DQ_RX_DATA_70to0[0] , LANE_0_IOD_DQ_RX_DATA_60to0[0] , LANE_0_IOD_DQ_RX_DATA_50to0[0] , LANE_0_IOD_DQ_RX_DATA_40to0[0] , LANE_0_IOD_DQ_RX_DATA_30to0[0] , LANE_0_IOD_DQ_RX_DATA_20to0[0] , LANE_0_IOD_DQ_RX_DATA_10to0[0] , LANE_0_IOD_DQ_RX_DATA_00to0[0] };
assign IOG_RDDATA_VALID_net_0          = { LANE_3_CTRL_RX_DATA_VALID , LANE_2_CTRL_RX_DATA_VALID , LANE_1_CTRL_RX_DATA_VALID , LANE_0_CTRL_RX_DATA_VALID };
assign PAD_RDDATA_net_0                = { LANE_3_IOD_DQ_RX_BYPASS_DATA_7 , LANE_3_IOD_DQ_RX_BYPASS_DATA_6 , LANE_3_IOD_DQ_RX_BYPASS_DATA_5 , LANE_3_IOD_DQ_RX_BYPASS_DATA_4 , LANE_3_IOD_DQ_RX_BYPASS_DATA_3 , LANE_3_IOD_DQ_RX_BYPASS_DATA_2 , LANE_3_IOD_DQ_RX_BYPASS_DATA_1 , LANE_3_IOD_DQ_RX_BYPASS_DATA_0 , LANE_2_IOD_DQ_RX_BYPASS_DATA_7 , LANE_2_IOD_DQ_RX_BYPASS_DATA_6 , LANE_2_IOD_DQ_RX_BYPASS_DATA_5 , LANE_2_IOD_DQ_RX_BYPASS_DATA_4 , LANE_2_IOD_DQ_RX_BYPASS_DATA_3 , LANE_2_IOD_DQ_RX_BYPASS_DATA_2 , LANE_2_IOD_DQ_RX_BYPASS_DATA_1 , LANE_2_IOD_DQ_RX_BYPASS_DATA_0 , LANE_1_IOD_DQ_RX_BYPASS_DATA_7 , LANE_1_IOD_DQ_RX_BYPASS_DATA_6 , LANE_1_IOD_DQ_RX_BYPASS_DATA_5 , LANE_1_IOD_DQ_RX_BYPASS_DATA_4 , LANE_1_IOD_DQ_RX_BYPASS_DATA_3 , LANE_1_IOD_DQ_RX_BYPASS_DATA_2 , LANE_1_IOD_DQ_RX_BYPASS_DATA_1 , LANE_1_IOD_DQ_RX_BYPASS_DATA_0 , LANE_0_IOD_DQ_RX_BYPASS_DATA_7 , LANE_0_IOD_DQ_RX_BYPASS_DATA_6 , LANE_0_IOD_DQ_RX_BYPASS_DATA_5 , LANE_0_IOD_DQ_RX_BYPASS_DATA_4 , LANE_0_IOD_DQ_RX_BYPASS_DATA_3 , LANE_0_IOD_DQ_RX_BYPASS_DATA_2 , LANE_0_IOD_DQ_RX_BYPASS_DATA_1 , LANE_0_IOD_DQ_RX_BYPASS_DATA_0 };
assign DQSW_EYE_MONITOR_EARLY_net_0    = { LANE_3_IOD_DQSW_TRAINING_EYE_MONITOR_EARLY_0 , LANE_2_IOD_DQSW_TRAINING_EYE_MONITOR_EARLY_0 , LANE_1_IOD_DQSW_TRAINING_EYE_MONITOR_EARLY_0 , LANE_0_IOD_DQSW_TRAINING_EYE_MONITOR_EARLY_0 };
assign DQSW_EYE_MONITOR_LATE_net_0     = { LANE_3_IOD_DQSW_TRAINING_EYE_MONITOR_LATE_0 , LANE_2_IOD_DQSW_TRAINING_EYE_MONITOR_LATE_0 , LANE_1_IOD_DQSW_TRAINING_EYE_MONITOR_LATE_0 , LANE_0_IOD_DQSW_TRAINING_EYE_MONITOR_LATE_0 };
assign DQSW270_EYE_MONITOR_EARLY_net_0 = { LANE_3_IOD_READ_TRAINING_EYE_MONITOR_EARLY_0 , LANE_2_IOD_READ_TRAINING_EYE_MONITOR_EARLY_0 , LANE_1_IOD_READ_TRAINING_EYE_MONITOR_EARLY_0 , LANE_0_IOD_READ_TRAINING_EYE_MONITOR_EARLY_0 };
assign DQSW270_EYE_MONITOR_LATE_net_0  = { LANE_3_IOD_READ_TRAINING_EYE_MONITOR_LATE_0 , LANE_2_IOD_READ_TRAINING_EYE_MONITOR_LATE_0 , LANE_1_IOD_READ_TRAINING_EYE_MONITOR_LATE_0 , LANE_0_IOD_READ_TRAINING_EYE_MONITOR_LATE_0 };
assign DQSW270_IGEAR_RX8_net_0         = { LANE_3_IOD_READ_TRAINING_RX_DATA_06to6[6] , LANE_2_IOD_READ_TRAINING_RX_DATA_06to6[6] , LANE_1_IOD_READ_TRAINING_RX_DATA_06to6[6] , LANE_0_IOD_READ_TRAINING_RX_DATA_06to6[6] };
assign DQSW_DELAY_LINE_OOR_net_0       = { LANE_3_IOD_DQSW_TRAINING_DELAY_LINE_OUT_OF_RANGE_0 , LANE_2_IOD_DQSW_TRAINING_DELAY_LINE_OUT_OF_RANGE_0 , LANE_1_IOD_DQSW_TRAINING_DELAY_LINE_OUT_OF_RANGE_0 , LANE_0_IOD_DQSW_TRAINING_DELAY_LINE_OUT_OF_RANGE_0 };
assign DQSW270_DELAY_LINE_OOR_net_0    = { LANE_3_IOD_READ_TRAINING_DELAY_LINE_OUT_OF_RANGE_0 , LANE_2_IOD_READ_TRAINING_DELAY_LINE_OUT_OF_RANGE_0 , LANE_1_IOD_READ_TRAINING_DELAY_LINE_OUT_OF_RANGE_0 , LANE_0_IOD_READ_TRAINING_DELAY_LINE_OUT_OF_RANGE_0 };
wire   [0:0]                               DFI_ADDRESS_P0_1919_unconnected;
wire   [0:0]                               DFI_ADDRESS_P0_1818_unconnected;
wire   [0:0]                               DFI_ADDRESS_P0_1717_unconnected;
wire   [0:0]                               DFI_ADDRESS_P0_1616_unconnected;
wire   [0:0]                               DFI_ADDRESS_P0_1515_unconnected;
wire   [0:0]                               DFI_ADDRESS_P0_1414_unconnected;
assign DFI_ADDRESS_P0_net_0            = { DFI_ADDRESS_P0_1919_unconnected , DFI_ADDRESS_P0_1818_unconnected , DFI_ADDRESS_P0_1717_unconnected , DFI_ADDRESS_P0_1616_unconnected , DFI_ADDRESS_P0_1515_unconnected , DFI_ADDRESS_P0_1414_unconnected , DFI_ADDRESS_P0_slice_13[13] , DFI_ADDRESS_P0_slice_12[12] , DFI_ADDRESS_P0_slice_11[11] , DFI_ADDRESS_P0_slice_10[10] , DFI_ADDRESS_P0_slice_9[9] , DFI_ADDRESS_P0_slice_8[8] , DFI_ADDRESS_P0_slice_7[7] , DFI_ADDRESS_P0_slice_6[6] , DFI_ADDRESS_P0_slice_5[5] , DFI_ADDRESS_P0_slice_4[4] , DFI_ADDRESS_P0_slice_3[3] , DFI_ADDRESS_P0_slice_2[2] , DFI_ADDRESS_P0_slice_1[1] , DFI_ADDRESS_P0_slice_0[0] };
wire   [0:0]                               DFI_ADDRESS_P1_1919_unconnected;
wire   [0:0]                               DFI_ADDRESS_P1_1818_unconnected;
wire   [0:0]                               DFI_ADDRESS_P1_1717_unconnected;
wire   [0:0]                               DFI_ADDRESS_P1_1616_unconnected;
wire   [0:0]                               DFI_ADDRESS_P1_1515_unconnected;
wire   [0:0]                               DFI_ADDRESS_P1_1414_unconnected;
assign DFI_ADDRESS_P1_net_0            = { DFI_ADDRESS_P1_1919_unconnected , DFI_ADDRESS_P1_1818_unconnected , DFI_ADDRESS_P1_1717_unconnected , DFI_ADDRESS_P1_1616_unconnected , DFI_ADDRESS_P1_1515_unconnected , DFI_ADDRESS_P1_1414_unconnected , DFI_ADDRESS_P1_slice_13[13] , DFI_ADDRESS_P1_slice_12[12] , DFI_ADDRESS_P1_slice_11[11] , DFI_ADDRESS_P1_slice_10[10] , DFI_ADDRESS_P1_slice_9[9] , DFI_ADDRESS_P1_slice_8[8] , DFI_ADDRESS_P1_slice_7[7] , DFI_ADDRESS_P1_slice_6[6] , DFI_ADDRESS_P1_slice_5[5] , DFI_ADDRESS_P1_slice_4[4] , DFI_ADDRESS_P1_slice_3[3] , DFI_ADDRESS_P1_slice_2[2] , DFI_ADDRESS_P1_slice_1[1] , DFI_ADDRESS_P1_slice_0[0] };
wire   [0:0]                               DFI_ADDRESS_P2_1919_unconnected;
wire   [0:0]                               DFI_ADDRESS_P2_1818_unconnected;
wire   [0:0]                               DFI_ADDRESS_P2_1717_unconnected;
wire   [0:0]                               DFI_ADDRESS_P2_1616_unconnected;
wire   [0:0]                               DFI_ADDRESS_P2_1515_unconnected;
wire   [0:0]                               DFI_ADDRESS_P2_1414_unconnected;
assign DFI_ADDRESS_P2_net_0            = { DFI_ADDRESS_P2_1919_unconnected , DFI_ADDRESS_P2_1818_unconnected , DFI_ADDRESS_P2_1717_unconnected , DFI_ADDRESS_P2_1616_unconnected , DFI_ADDRESS_P2_1515_unconnected , DFI_ADDRESS_P2_1414_unconnected , DFI_ADDRESS_P2_slice_13[13] , DFI_ADDRESS_P2_slice_12[12] , DFI_ADDRESS_P2_slice_11[11] , DFI_ADDRESS_P2_slice_10[10] , DFI_ADDRESS_P2_slice_9[9] , DFI_ADDRESS_P2_slice_8[8] , DFI_ADDRESS_P2_slice_7[7] , DFI_ADDRESS_P2_slice_6[6] , DFI_ADDRESS_P2_slice_5[5] , DFI_ADDRESS_P2_slice_4[4] , DFI_ADDRESS_P2_slice_3[3] , DFI_ADDRESS_P2_slice_2[2] , DFI_ADDRESS_P2_slice_1[1] , DFI_ADDRESS_P2_slice_0[0] };
wire   [0:0]                               DFI_ADDRESS_P3_1919_unconnected;
wire   [0:0]                               DFI_ADDRESS_P3_1818_unconnected;
wire   [0:0]                               DFI_ADDRESS_P3_1717_unconnected;
wire   [0:0]                               DFI_ADDRESS_P3_1616_unconnected;
wire   [0:0]                               DFI_ADDRESS_P3_1515_unconnected;
wire   [0:0]                               DFI_ADDRESS_P3_1414_unconnected;
assign DFI_ADDRESS_P3_net_0            = { DFI_ADDRESS_P3_1919_unconnected , DFI_ADDRESS_P3_1818_unconnected , DFI_ADDRESS_P3_1717_unconnected , DFI_ADDRESS_P3_1616_unconnected , DFI_ADDRESS_P3_1515_unconnected , DFI_ADDRESS_P3_1414_unconnected , DFI_ADDRESS_P3_slice_13[13] , DFI_ADDRESS_P3_slice_12[12] , DFI_ADDRESS_P3_slice_11[11] , DFI_ADDRESS_P3_slice_10[10] , DFI_ADDRESS_P3_slice_9[9] , DFI_ADDRESS_P3_slice_8[8] , DFI_ADDRESS_P3_slice_7[7] , DFI_ADDRESS_P3_slice_6[6] , DFI_ADDRESS_P3_slice_5[5] , DFI_ADDRESS_P3_slice_4[4] , DFI_ADDRESS_P3_slice_3[3] , DFI_ADDRESS_P3_slice_2[2] , DFI_ADDRESS_P3_slice_1[1] , DFI_ADDRESS_P3_slice_0[0] };
assign BCLK_IGEAR_RX_net_0             = { IOD_BCLK_TRAINING_RX_DATA_06to6[6] , IOD_BCLK_TRAINING_RX_DATA_04to4[4] , IOD_BCLK_TRAINING_RX_DATA_02to2[2] , IOD_BCLK_TRAINING_RX_DATA_00to0[0] };
assign DQSW270_IGEAR_RX_net_0          = { LANE_3_IOD_READ_TRAINING_RX_DATA_07to7[7] , LANE_3_IOD_READ_TRAINING_RX_DATA_06to6[6] , LANE_2_IOD_READ_TRAINING_RX_DATA_07to7[7] , LANE_2_IOD_READ_TRAINING_RX_DATA_06to6[6] , LANE_1_IOD_READ_TRAINING_RX_DATA_07to7[7] , LANE_1_IOD_READ_TRAINING_RX_DATA_06to6[6] , LANE_0_IOD_READ_TRAINING_RX_DATA_07to7[7] , LANE_0_IOD_READ_TRAINING_RX_DATA_06to6[6] };
assign DQSW_IGEAR_RX_net_0             = { LANE_3_IOD_DQSW_TRAINING_RX_DATA_01to1[1] , LANE_3_IOD_DQSW_TRAINING_RX_DATA_00to0[0] , LANE_2_IOD_DQSW_TRAINING_RX_DATA_01to1[1] , LANE_2_IOD_DQSW_TRAINING_RX_DATA_00to0[0] , LANE_1_IOD_DQSW_TRAINING_RX_DATA_01to1[1] , LANE_1_IOD_DQSW_TRAINING_RX_DATA_00to0[0] , LANE_0_IOD_DQSW_TRAINING_RX_DATA_01to1[1] , LANE_0_IOD_DQSW_TRAINING_RX_DATA_00to0[0] };
assign IOG_DQ_TXDATA_IN_net_0          = { DFI_WRDATA_P3_slice_63[63] , DFI_WRDATA_P3_slice_62[31] , DFI_WRDATA_P2_slice_63[63] , DFI_WRDATA_P2_slice_62[31] , DFI_WRDATA_P1_slice_63[63] , DFI_WRDATA_P1_slice_62[31] , DFI_WRDATA_P0_slice_63[63] , DFI_WRDATA_P0_slice_62[31] , DFI_WRDATA_P3_slice_61[62] , DFI_WRDATA_P3_slice_60[30] , DFI_WRDATA_P2_slice_61[62] , DFI_WRDATA_P2_slice_60[30] , DFI_WRDATA_P1_slice_61[62] , DFI_WRDATA_P1_slice_60[30] , DFI_WRDATA_P0_slice_61[62] , DFI_WRDATA_P0_slice_60[30] , DFI_WRDATA_P3_slice_59[61] , DFI_WRDATA_P3_slice_58[29] , DFI_WRDATA_P2_slice_59[61] , DFI_WRDATA_P2_slice_58[29] , DFI_WRDATA_P1_slice_59[61] , DFI_WRDATA_P1_slice_58[29] , DFI_WRDATA_P0_slice_59[61] , DFI_WRDATA_P0_slice_58[29] , DFI_WRDATA_P3_slice_57[60] , DFI_WRDATA_P3_slice_56[28] , DFI_WRDATA_P2_slice_57[60] , DFI_WRDATA_P2_slice_56[28] , DFI_WRDATA_P1_slice_57[60] , DFI_WRDATA_P1_slice_56[28] , DFI_WRDATA_P0_slice_57[60] , DFI_WRDATA_P0_slice_56[28] , DFI_WRDATA_P3_slice_55[59] , DFI_WRDATA_P3_slice_54[27] , DFI_WRDATA_P2_slice_55[59] , DFI_WRDATA_P2_slice_54[27] , DFI_WRDATA_P1_slice_55[59] , DFI_WRDATA_P1_slice_54[27] , DFI_WRDATA_P0_slice_55[59] , DFI_WRDATA_P0_slice_54[27] , DFI_WRDATA_P3_slice_53[58] , DFI_WRDATA_P3_slice_52[26] , DFI_WRDATA_P2_slice_53[58] , DFI_WRDATA_P2_slice_52[26] , DFI_WRDATA_P1_slice_53[58] , DFI_WRDATA_P1_slice_52[26] , DFI_WRDATA_P0_slice_53[58] , DFI_WRDATA_P0_slice_52[26] , DFI_WRDATA_P3_slice_51[57] , DFI_WRDATA_P3_slice_50[25] , DFI_WRDATA_P2_slice_51[57] , DFI_WRDATA_P2_slice_50[25] , DFI_WRDATA_P1_slice_51[57] , DFI_WRDATA_P1_slice_50[25] , DFI_WRDATA_P0_slice_51[57] , DFI_WRDATA_P0_slice_50[25] , DFI_WRDATA_P3_slice_49[56] , DFI_WRDATA_P3_slice_48[24] , DFI_WRDATA_P2_slice_49[56] , DFI_WRDATA_P2_slice_48[24] , DFI_WRDATA_P1_slice_49[56] , DFI_WRDATA_P1_slice_48[24] , DFI_WRDATA_P0_slice_49[56] , DFI_WRDATA_P0_slice_48[24] , DFI_WRDATA_P3_slice_47[55] , DFI_WRDATA_P3_slice_46[23] , DFI_WRDATA_P2_slice_47[55] , DFI_WRDATA_P2_slice_46[23] , DFI_WRDATA_P1_slice_47[55] , DFI_WRDATA_P1_slice_46[23] , DFI_WRDATA_P0_slice_47[55] , DFI_WRDATA_P0_slice_46[23] , DFI_WRDATA_P3_slice_45[54] , DFI_WRDATA_P3_slice_44[22] , DFI_WRDATA_P2_slice_45[54] , DFI_WRDATA_P2_slice_44[22] , DFI_WRDATA_P1_slice_45[54] , DFI_WRDATA_P1_slice_44[22] , DFI_WRDATA_P0_slice_45[54] , DFI_WRDATA_P0_slice_44[22] , DFI_WRDATA_P3_slice_43[53] , DFI_WRDATA_P3_slice_42[21] , DFI_WRDATA_P2_slice_43[53] , DFI_WRDATA_P2_slice_42[21] , DFI_WRDATA_P1_slice_43[53] , DFI_WRDATA_P1_slice_42[21] , DFI_WRDATA_P0_slice_43[53] , DFI_WRDATA_P0_slice_42[21] , DFI_WRDATA_P3_slice_41[52] , DFI_WRDATA_P3_slice_40[20] , DFI_WRDATA_P2_slice_41[52] , DFI_WRDATA_P2_slice_40[20] , DFI_WRDATA_P1_slice_41[52] , DFI_WRDATA_P1_slice_40[20] , DFI_WRDATA_P0_slice_41[52] , DFI_WRDATA_P0_slice_40[20] , DFI_WRDATA_P3_slice_39[51] , DFI_WRDATA_P3_slice_38[19] , DFI_WRDATA_P2_slice_39[51] , DFI_WRDATA_P2_slice_38[19] , DFI_WRDATA_P1_slice_39[51] , DFI_WRDATA_P1_slice_38[19] , DFI_WRDATA_P0_slice_39[51] , DFI_WRDATA_P0_slice_38[19] , DFI_WRDATA_P3_slice_37[50] , DFI_WRDATA_P3_slice_36[18] , DFI_WRDATA_P2_slice_37[50] , DFI_WRDATA_P2_slice_36[18] , DFI_WRDATA_P1_slice_37[50] , DFI_WRDATA_P1_slice_36[18] , DFI_WRDATA_P0_slice_37[50] , DFI_WRDATA_P0_slice_36[18] , DFI_WRDATA_P3_slice_35[49] , DFI_WRDATA_P3_slice_34[17] , DFI_WRDATA_P2_slice_35[49] , DFI_WRDATA_P2_slice_34[17] , DFI_WRDATA_P1_slice_35[49] , DFI_WRDATA_P1_slice_34[17] , DFI_WRDATA_P0_slice_35[49] , DFI_WRDATA_P0_slice_34[17] , DFI_WRDATA_P3_slice_33[48] , DFI_WRDATA_P3_slice_32[16] , DFI_WRDATA_P2_slice_33[48] , DFI_WRDATA_P2_slice_32[16] , DFI_WRDATA_P1_slice_33[48] , DFI_WRDATA_P1_slice_32[16] , DFI_WRDATA_P0_slice_33[48] , DFI_WRDATA_P0_slice_32[16] , DFI_WRDATA_P3_slice_31[47] , DFI_WRDATA_P3_slice_30[15] , DFI_WRDATA_P2_slice_31[47] , DFI_WRDATA_P2_slice_30[15] , DFI_WRDATA_P1_slice_31[47] , DFI_WRDATA_P1_slice_30[15] , DFI_WRDATA_P0_slice_31[47] , DFI_WRDATA_P0_slice_30[15] , DFI_WRDATA_P3_slice_29[46] , DFI_WRDATA_P3_slice_28[14] , DFI_WRDATA_P2_slice_29[46] , DFI_WRDATA_P2_slice_28[14] , DFI_WRDATA_P1_slice_29[46] , DFI_WRDATA_P1_slice_28[14] , DFI_WRDATA_P0_slice_29[46] , DFI_WRDATA_P0_slice_28[14] , DFI_WRDATA_P3_slice_27[45] , DFI_WRDATA_P3_slice_26[13] , DFI_WRDATA_P2_slice_27[45] , DFI_WRDATA_P2_slice_26[13] , DFI_WRDATA_P1_slice_27[45] , DFI_WRDATA_P1_slice_26[13] , DFI_WRDATA_P0_slice_27[45] , DFI_WRDATA_P0_slice_26[13] , DFI_WRDATA_P3_slice_25[44] , DFI_WRDATA_P3_slice_24[12] , DFI_WRDATA_P2_slice_25[44] , DFI_WRDATA_P2_slice_24[12] , DFI_WRDATA_P1_slice_25[44] , DFI_WRDATA_P1_slice_24[12] , DFI_WRDATA_P0_slice_25[44] , DFI_WRDATA_P0_slice_24[12] , DFI_WRDATA_P3_slice_23[43] , DFI_WRDATA_P3_slice_22[11] , DFI_WRDATA_P2_slice_23[43] , DFI_WRDATA_P2_slice_22[11] , DFI_WRDATA_P1_slice_23[43] , DFI_WRDATA_P1_slice_22[11] , DFI_WRDATA_P0_slice_23[43] , DFI_WRDATA_P0_slice_22[11] , DFI_WRDATA_P3_slice_21[42] , DFI_WRDATA_P3_slice_20[10] , DFI_WRDATA_P2_slice_21[42] , DFI_WRDATA_P2_slice_20[10] , DFI_WRDATA_P1_slice_21[42] , DFI_WRDATA_P1_slice_20[10] , DFI_WRDATA_P0_slice_21[42] , DFI_WRDATA_P0_slice_20[10] , DFI_WRDATA_P3_slice_19[41] , DFI_WRDATA_P3_slice_18[9] , DFI_WRDATA_P2_slice_19[41] , DFI_WRDATA_P2_slice_18[9] , DFI_WRDATA_P1_slice_19[41] , DFI_WRDATA_P1_slice_18[9] , DFI_WRDATA_P0_slice_19[41] , DFI_WRDATA_P0_slice_18[9] , DFI_WRDATA_P3_slice_17[40] , DFI_WRDATA_P3_slice_16[8] , DFI_WRDATA_P2_slice_17[40] , DFI_WRDATA_P2_slice_16[8] , DFI_WRDATA_P1_slice_17[40] , DFI_WRDATA_P1_slice_16[8] , DFI_WRDATA_P0_slice_17[40] , DFI_WRDATA_P0_slice_16[8] , DFI_WRDATA_P3_slice_15[39] , DFI_WRDATA_P3_slice_14[7] , DFI_WRDATA_P2_slice_15[39] , DFI_WRDATA_P2_slice_14[7] , DFI_WRDATA_P1_slice_15[39] , DFI_WRDATA_P1_slice_14[7] , DFI_WRDATA_P0_slice_15[39] , DFI_WRDATA_P0_slice_14[7] , DFI_WRDATA_P3_slice_13[38] , DFI_WRDATA_P3_slice_12[6] , DFI_WRDATA_P2_slice_13[38] , DFI_WRDATA_P2_slice_12[6] , DFI_WRDATA_P1_slice_13[38] , DFI_WRDATA_P1_slice_12[6] , DFI_WRDATA_P0_slice_13[38] , DFI_WRDATA_P0_slice_12[6] , DFI_WRDATA_P3_slice_11[37] , DFI_WRDATA_P3_slice_10[5] , DFI_WRDATA_P2_slice_11[37] , DFI_WRDATA_P2_slice_10[5] , DFI_WRDATA_P1_slice_11[37] , DFI_WRDATA_P1_slice_10[5] , DFI_WRDATA_P0_slice_11[37] , DFI_WRDATA_P0_slice_10[5] , DFI_WRDATA_P3_slice_9[36] , DFI_WRDATA_P3_slice_8[4] , DFI_WRDATA_P2_slice_9[36] , DFI_WRDATA_P2_slice_8[4] , DFI_WRDATA_P1_slice_9[36] , DFI_WRDATA_P1_slice_8[4] , DFI_WRDATA_P0_slice_9[36] , DFI_WRDATA_P0_slice_8[4] , DFI_WRDATA_P3_slice_7[35] , DFI_WRDATA_P3_slice_6[3] , DFI_WRDATA_P2_slice_7[35] , DFI_WRDATA_P2_slice_6[3] , DFI_WRDATA_P1_slice_7[35] , DFI_WRDATA_P1_slice_6[3] , DFI_WRDATA_P0_slice_7[35] , DFI_WRDATA_P0_slice_6[3] , DFI_WRDATA_P3_slice_5[34] , DFI_WRDATA_P3_slice_4[2] , DFI_WRDATA_P2_slice_5[34] , DFI_WRDATA_P2_slice_4[2] , DFI_WRDATA_P1_slice_5[34] , DFI_WRDATA_P1_slice_4[2] , DFI_WRDATA_P0_slice_5[34] , DFI_WRDATA_P0_slice_4[2] , DFI_WRDATA_P3_slice_3[33] , DFI_WRDATA_P3_slice_2[1] , DFI_WRDATA_P2_slice_3[33] , DFI_WRDATA_P2_slice_2[1] , DFI_WRDATA_P1_slice_3[33] , DFI_WRDATA_P1_slice_2[1] , DFI_WRDATA_P0_slice_3[33] , DFI_WRDATA_P0_slice_2[1] , DFI_WRDATA_P3_slice_1[32] , DFI_WRDATA_P3_slice_0[0] , DFI_WRDATA_P2_slice_1[32] , DFI_WRDATA_P2_slice_0[0] , DFI_WRDATA_P1_slice_1[32] , DFI_WRDATA_P1_slice_0[0] , DFI_WRDATA_P0_slice_1[32] , DFI_WRDATA_P0_slice_0[0] };
assign IOG_DM_TXDATA_IN_net_0          = { DFI_WRDATA_MASK_P3_slice_7[7] , DFI_WRDATA_MASK_P3_slice_6[3] , DFI_WRDATA_MASK_P2_slice_7[7] , DFI_WRDATA_MASK_P2_slice_6[3] , DFI_WRDATA_MASK_P1_slice_7[7] , DFI_WRDATA_MASK_P1_slice_6[3] , DFI_WRDATA_MASK_P0_slice_7[7] , DFI_WRDATA_MASK_P0_slice_6[3] , DFI_WRDATA_MASK_P3_slice_5[6] , DFI_WRDATA_MASK_P3_slice_4[2] , DFI_WRDATA_MASK_P2_slice_5[6] , DFI_WRDATA_MASK_P2_slice_4[2] , DFI_WRDATA_MASK_P1_slice_5[6] , DFI_WRDATA_MASK_P1_slice_4[2] , DFI_WRDATA_MASK_P0_slice_5[6] , DFI_WRDATA_MASK_P0_slice_4[2] , DFI_WRDATA_MASK_P3_slice_3[5] , DFI_WRDATA_MASK_P3_slice_2[1] , DFI_WRDATA_MASK_P2_slice_3[5] , DFI_WRDATA_MASK_P2_slice_2[1] , DFI_WRDATA_MASK_P1_slice_3[5] , DFI_WRDATA_MASK_P1_slice_2[1] , DFI_WRDATA_MASK_P0_slice_3[5] , DFI_WRDATA_MASK_P0_slice_2[1] , DFI_WRDATA_MASK_P3_slice_1[4] , DFI_WRDATA_MASK_P3_slice_0[0] , DFI_WRDATA_MASK_P2_slice_1[4] , DFI_WRDATA_MASK_P2_slice_0[0] , DFI_WRDATA_MASK_P1_slice_1[4] , DFI_WRDATA_MASK_P1_slice_0[0] , DFI_WRDATA_MASK_P0_slice_1[4] , DFI_WRDATA_MASK_P0_slice_0[0] };
wire   [0:0]                          DFI_BANK_P0_22_unconnected;
assign DFI_BANK_P0_net_0               = { DFI_BANK_P0_22_unconnected , DFI_BANK_P0_slice_1[1] , DFI_BANK_P0_slice_0[0] };
wire   [0:0]                          DFI_BANK_P1_22_unconnected;
assign DFI_BANK_P1_net_0               = { DFI_BANK_P1_22_unconnected , DFI_BANK_P1_slice_1[1] , DFI_BANK_P1_slice_0[0] };
wire   [0:0]                          DFI_BANK_P2_22_unconnected;
assign DFI_BANK_P2_net_0               = { DFI_BANK_P2_22_unconnected , DFI_BANK_P2_slice_1[1] , DFI_BANK_P2_slice_0[0] };
wire   [0:0]                          DFI_BANK_P3_22_unconnected;
assign DFI_BANK_P3_net_0               = { DFI_BANK_P3_22_unconnected , DFI_BANK_P3_slice_1[1] , DFI_BANK_P3_slice_0[0] };
assign DFI_BG_P0_net_0                 = { DFI_BG_P0_slice_1[1] , DFI_BG_P0_slice_0[0] };
assign DFI_BG_P1_net_0                 = { DFI_BG_P1_slice_1[1] , DFI_BG_P1_slice_0[0] };
assign DFI_BG_P2_net_0                 = { DFI_BG_P2_slice_1[1] , DFI_BG_P2_slice_0[0] };
assign DFI_BG_P3_net_0                 = { DFI_BG_P3_slice_1[1] , DFI_BG_P3_slice_0[0] };
assign PAD_net_0                       = { DQ[7:7] , DQ[6:6] , DQ[5:5] , DQ[4:4] , DQ[3:3] , DQ[2:2] , DQ[1:1] , DQ[0:0] };
assign PAD_net_1                       = { DQ[15:15] , DQ[14:14] , DQ[13:13] , DQ[12:12] , DQ[11:11] , DQ[10:10] , DQ[9:9] , DQ[8:8] };
assign PAD_net_2                       = { DQ[23:23] , DQ[22:22] , DQ[21:21] , DQ[20:20] , DQ[19:19] , DQ[18:18] , DQ[17:17] , DQ[16:16] };
assign PAD_net_3                       = { DQ[31:31] , DQ[30:30] , DQ[29:29] , DQ[28:28] , DQ[27:27] , DQ[26:26] , DQ[25:25] , DQ[24:24] };
//--------------------------------------------------------------------
// Component instances
//--------------------------------------------------------------------
//--------CLKINT_PRESERVE
CLKINT_PRESERVE CLKINT_CMD(
        // Inputs
        .A ( DFN1_CMD_Q ),
        // Outputs
        .Y ( CLKINT_CMD_Y ) 
        );

//--------DFN1
DFN1 DFN1_CMD(
        // Inputs
        .D   ( IOD_TRAINING_0_CMD_RESET_LANE ),
        .CLK ( SYS_CLK ),
        // Outputs
        .Q   ( DFN1_CMD_Q ) 
        );

//--------PF_DDR4_SS_DDRPHY_BLK_IOD_A_11_0_PF_IOD   -   Actel:SgCore:PF_IOD:1.0.218
PF_DDR4_SS_DDRPHY_BLK_IOD_A_11_0_PF_IOD IOD_A_11_0(
        // Inputs
        .ARST_N                     ( LANECTRL_ADDR_CMD_0_ARST_N ),
        .RX_SYNC_RST                ( LANECTRL_ADDR_CMD_0_RX_SYNC_RST ),
        .TX_SYNC_RST                ( LANECTRL_ADDR_CMD_0_TX_SYNC_RST ),
        .HS_IO_CLK                  ( HS_IO_CLK ),
        .TX_DQS_270                 ( LANECTRL_ADDR_CMD_0_TX_DQS_270 ),
        .TX_DATA_0                  ( TX_DATA_0_net_0 ),
        .TX_DATA_1                  ( TX_DATA_1_net_0 ),
        .TX_DATA_2                  ( TX_DATA_2_net_0 ),
        .TX_DATA_3                  ( TX_DATA_3_net_0 ),
        .TX_DATA_4                  ( TX_DATA_4_net_0 ),
        .TX_DATA_5                  ( TX_DATA_5_net_0 ),
        .TX_DATA_6                  ( TX_DATA_6_net_0 ),
        .TX_DATA_7                  ( TX_DATA_7_net_0 ),
        .TX_DATA_8                  ( TX_DATA_8_net_0 ),
        .TX_DATA_9                  ( TX_DATA_9_net_0 ),
        .TX_DATA_10                 ( TX_DATA_10_net_0 ),
        .TX_DATA_11                 ( TX_DATA_11_net_0 ),
        .OE_DATA_0                  ( OE_DATA_0_const_net_0 ),
        .OE_DATA_1                  ( OE_DATA_1_const_net_0 ),
        .OE_DATA_2                  ( OE_DATA_2_const_net_0 ),
        .OE_DATA_3                  ( OE_DATA_3_const_net_0 ),
        .OE_DATA_4                  ( OE_DATA_4_const_net_0 ),
        .OE_DATA_5                  ( OE_DATA_5_const_net_0 ),
        .OE_DATA_6                  ( OE_DATA_6_const_net_0 ),
        .OE_DATA_7                  ( OE_DATA_7_const_net_0 ),
        .OE_DATA_8                  ( OE_DATA_8_const_net_0 ),
        .OE_DATA_9                  ( OE_DATA_9_const_net_0 ),
        .OE_DATA_10                 ( OE_DATA_10_const_net_0 ),
        .OE_DATA_11                 ( OE_DATA_11_const_net_0 ),
        .DELAY_LINE_MOVE_0          ( IOD_TRAINING_0_CMD_DELAY_LINE_MOVE ),
        .DELAY_LINE_MOVE_1          ( IOD_TRAINING_0_CMD_DELAY_LINE_MOVE ),
        .DELAY_LINE_MOVE_2          ( IOD_TRAINING_0_CMD_DELAY_LINE_MOVE ),
        .DELAY_LINE_MOVE_3          ( IOD_TRAINING_0_CMD_DELAY_LINE_MOVE ),
        .DELAY_LINE_MOVE_4          ( IOD_TRAINING_0_CMD_DELAY_LINE_MOVE ),
        .DELAY_LINE_MOVE_5          ( IOD_TRAINING_0_CMD_DELAY_LINE_MOVE ),
        .DELAY_LINE_MOVE_6          ( IOD_TRAINING_0_CMD_DELAY_LINE_MOVE ),
        .DELAY_LINE_MOVE_7          ( IOD_TRAINING_0_CMD_DELAY_LINE_MOVE ),
        .DELAY_LINE_MOVE_8          ( IOD_TRAINING_0_CMD_DELAY_LINE_MOVE ),
        .DELAY_LINE_MOVE_9          ( IOD_TRAINING_0_CMD_DELAY_LINE_MOVE ),
        .DELAY_LINE_MOVE_10         ( IOD_TRAINING_0_CMD_DELAY_LINE_MOVE ),
        .DELAY_LINE_MOVE_11         ( IOD_TRAINING_0_CMD_DELAY_LINE_MOVE ),
        .DELAY_LINE_DIRECTION_0     ( IOD_TRAINING_0_CMD_DELAY_LINE_DIRECTION ),
        .DELAY_LINE_DIRECTION_1     ( IOD_TRAINING_0_CMD_DELAY_LINE_DIRECTION ),
        .DELAY_LINE_DIRECTION_2     ( IOD_TRAINING_0_CMD_DELAY_LINE_DIRECTION ),
        .DELAY_LINE_DIRECTION_3     ( IOD_TRAINING_0_CMD_DELAY_LINE_DIRECTION ),
        .DELAY_LINE_DIRECTION_4     ( IOD_TRAINING_0_CMD_DELAY_LINE_DIRECTION ),
        .DELAY_LINE_DIRECTION_5     ( IOD_TRAINING_0_CMD_DELAY_LINE_DIRECTION ),
        .DELAY_LINE_DIRECTION_6     ( IOD_TRAINING_0_CMD_DELAY_LINE_DIRECTION ),
        .DELAY_LINE_DIRECTION_7     ( IOD_TRAINING_0_CMD_DELAY_LINE_DIRECTION ),
        .DELAY_LINE_DIRECTION_8     ( IOD_TRAINING_0_CMD_DELAY_LINE_DIRECTION ),
        .DELAY_LINE_DIRECTION_9     ( IOD_TRAINING_0_CMD_DELAY_LINE_DIRECTION ),
        .DELAY_LINE_DIRECTION_10    ( IOD_TRAINING_0_CMD_DELAY_LINE_DIRECTION ),
        .DELAY_LINE_DIRECTION_11    ( IOD_TRAINING_0_CMD_DELAY_LINE_DIRECTION ),
        .DELAY_LINE_LOAD_0          ( IOD_TRAINING_0_CMD_DELAY_LINE_LOAD ),
        .DELAY_LINE_LOAD_1          ( IOD_TRAINING_0_CMD_DELAY_LINE_LOAD ),
        .DELAY_LINE_LOAD_2          ( IOD_TRAINING_0_CMD_DELAY_LINE_LOAD ),
        .DELAY_LINE_LOAD_3          ( IOD_TRAINING_0_CMD_DELAY_LINE_LOAD ),
        .DELAY_LINE_LOAD_4          ( IOD_TRAINING_0_CMD_DELAY_LINE_LOAD ),
        .DELAY_LINE_LOAD_5          ( IOD_TRAINING_0_CMD_DELAY_LINE_LOAD ),
        .DELAY_LINE_LOAD_6          ( IOD_TRAINING_0_CMD_DELAY_LINE_LOAD ),
        .DELAY_LINE_LOAD_7          ( IOD_TRAINING_0_CMD_DELAY_LINE_LOAD ),
        .DELAY_LINE_LOAD_8          ( IOD_TRAINING_0_CMD_DELAY_LINE_LOAD ),
        .DELAY_LINE_LOAD_9          ( IOD_TRAINING_0_CMD_DELAY_LINE_LOAD ),
        .DELAY_LINE_LOAD_10         ( IOD_TRAINING_0_CMD_DELAY_LINE_LOAD ),
        .DELAY_LINE_LOAD_11         ( IOD_TRAINING_0_CMD_DELAY_LINE_LOAD ),
        .FAB_CLK                    ( SYS_CLK ),
        .ODT_EN_0                   ( GND_net ), // tied to 1'b0 from definition
        .ODT_EN_1                   ( GND_net ), // tied to 1'b0 from definition
        .ODT_EN_2                   ( GND_net ), // tied to 1'b0 from definition
        .ODT_EN_3                   ( GND_net ), // tied to 1'b0 from definition
        .ODT_EN_4                   ( GND_net ), // tied to 1'b0 from definition
        .ODT_EN_5                   ( GND_net ), // tied to 1'b0 from definition
        .ODT_EN_6                   ( GND_net ), // tied to 1'b0 from definition
        .ODT_EN_7                   ( GND_net ), // tied to 1'b0 from definition
        .ODT_EN_8                   ( GND_net ), // tied to 1'b0 from definition
        .ODT_EN_9                   ( GND_net ), // tied to 1'b0 from definition
        .ODT_EN_10                  ( GND_net ), // tied to 1'b0 from definition
        .ODT_EN_11                  ( GND_net ), // tied to 1'b0 from definition
        // Outputs
        .DELAY_LINE_OUT_OF_RANGE_0  (  ),
        .DELAY_LINE_OUT_OF_RANGE_1  (  ),
        .DELAY_LINE_OUT_OF_RANGE_2  (  ),
        .DELAY_LINE_OUT_OF_RANGE_3  (  ),
        .DELAY_LINE_OUT_OF_RANGE_4  (  ),
        .DELAY_LINE_OUT_OF_RANGE_5  (  ),
        .DELAY_LINE_OUT_OF_RANGE_6  (  ),
        .DELAY_LINE_OUT_OF_RANGE_7  (  ),
        .DELAY_LINE_OUT_OF_RANGE_8  (  ),
        .DELAY_LINE_OUT_OF_RANGE_9  (  ),
        .DELAY_LINE_OUT_OF_RANGE_10 (  ),
        .DELAY_LINE_OUT_OF_RANGE_11 (  ),
        .PAD_O                      ( PAD_O_net_0 ) 
        );

//--------PF_DDR4_SS_DDRPHY_BLK_IOD_A_12_PF_IOD   -   Actel:SgCore:PF_IOD:1.0.218
PF_DDR4_SS_DDRPHY_BLK_IOD_A_12_PF_IOD IOD_A_12(
        // Inputs
        .RX_P_0                    ( OB_A_12_Y ),
        .ARST_N                    ( LANECTRL_ADDR_CMD_0_ARST_N ),
        .RX_SYNC_RST               ( LANECTRL_ADDR_CMD_0_RX_SYNC_RST ),
        .TX_SYNC_RST               ( LANECTRL_ADDR_CMD_0_TX_SYNC_RST ),
        .HS_IO_CLK                 ( HS_IO_CLK ),
        .TX_DQS_270                ( LANECTRL_ADDR_CMD_0_TX_DQS_270 ),
        .TX_DATA_0                 ( TX_DATA_0_net_1 ),
        .OE_DATA_0                 ( OE_DATA_0_net_0 ),
        .EYE_MONITOR_CLEAR_FLAGS_0 ( IOD_TRAINING_0_CMD_EYE_MONITOR_CLR_FLAGS ),
        .DELAY_LINE_MOVE_0         ( IOD_TRAINING_0_CMD_DELAY_LINE_MOVE_TRN ),
        .DELAY_LINE_DIRECTION_0    ( IOD_TRAINING_0_CMD_DELAY_LINE_DIRECTION ),
        .DELAY_LINE_LOAD_0         ( IOD_TRAINING_0_CMD_DELAY_LINE_LOAD ),
        .FAB_CLK                   ( SYS_CLK ),
        .ODT_EN_0                  ( GND_net ), // tied to 1'b0 from definition
        // Outputs
        .TX_0                      ( IOD_A_12_TX_0 ),
        .OE_0                      (  ),
        .DELAY_LINE_OUT_OF_RANGE_0 (  ),
        .EYE_MONITOR_EARLY_0       ( IOD_A_12_EYE_MONITOR_EARLY_0 ),
        .EYE_MONITOR_LATE_0        ( IOD_A_12_EYE_MONITOR_LATE_0 ),
        .RX_DATA_0                 ( RX_DATA_0_net_0 ) 
        );

//--------PF_DDR4_SS_DDRPHY_BLK_IOD_A_13_PF_IOD   -   Actel:SgCore:PF_IOD:1.0.218
PF_DDR4_SS_DDRPHY_BLK_IOD_A_13_PF_IOD IOD_A_13(
        // Inputs
        .ARST_N                    ( LANECTRL_ADDR_CMD_0_ARST_N ),
        .RX_SYNC_RST               ( LANECTRL_ADDR_CMD_0_RX_SYNC_RST ),
        .TX_SYNC_RST               ( LANECTRL_ADDR_CMD_0_TX_SYNC_RST ),
        .HS_IO_CLK                 ( HS_IO_CLK ),
        .TX_DQS_270                ( LANECTRL_ADDR_CMD_0_TX_DQS_270 ),
        .TX_DATA_0                 ( TX_DATA_0_net_2 ),
        .OE_DATA_0                 ( OE_DATA_0_const_net_1 ),
        .DELAY_LINE_MOVE_0         ( IOD_TRAINING_0_CMD_DELAY_LINE_MOVE ),
        .DELAY_LINE_DIRECTION_0    ( IOD_TRAINING_0_CMD_DELAY_LINE_DIRECTION ),
        .DELAY_LINE_LOAD_0         ( IOD_TRAINING_0_CMD_DELAY_LINE_LOAD ),
        .FAB_CLK                   ( SYS_CLK ),
        .ODT_EN_0                  ( GND_net ), // tied to 1'b0 from definition
        // Outputs
        .DELAY_LINE_OUT_OF_RANGE_0 (  ),
        .PAD_O                     ( A_12 ) 
        );

//--------PF_DDR4_SS_DDRPHY_BLK_IOD_ACT_N_PF_IOD   -   Actel:SgCore:PF_IOD:1.0.218
PF_DDR4_SS_DDRPHY_BLK_IOD_ACT_N_PF_IOD IOD_ACT_N(
        // Inputs
        .ARST_N                    ( LANECTRL_ADDR_CMD_0_ARST_N ),
        .RX_SYNC_RST               ( LANECTRL_ADDR_CMD_0_RX_SYNC_RST ),
        .TX_SYNC_RST               ( LANECTRL_ADDR_CMD_0_TX_SYNC_RST ),
        .HS_IO_CLK                 ( HS_IO_CLK ),
        .TX_DQS_270                ( LANECTRL_ADDR_CMD_0_TX_DQS_270 ),
        .TX_DATA_0                 ( TX_DATA_0_net_3 ),
        .OE_DATA_0                 ( OE_DATA_0_const_net_2 ),
        .DELAY_LINE_MOVE_0         ( IOD_TRAINING_0_CMD_DELAY_LINE_MOVE ),
        .DELAY_LINE_DIRECTION_0    ( IOD_TRAINING_0_CMD_DELAY_LINE_DIRECTION ),
        .DELAY_LINE_LOAD_0         ( IOD_TRAINING_0_CMD_DELAY_LINE_LOAD ),
        .FAB_CLK                   ( SYS_CLK ),
        .ODT_EN_0                  ( GND_net ), // tied to 1'b0 from definition
        // Outputs
        .DELAY_LINE_OUT_OF_RANGE_0 (  ),
        .PAD_O                     ( ACT_N_net_0 ) 
        );

//--------PF_DDR4_SS_DDRPHY_BLK_IOD_BA_PF_IOD   -   Actel:SgCore:PF_IOD:1.0.218
PF_DDR4_SS_DDRPHY_BLK_IOD_BA_PF_IOD IOD_BA(
        // Inputs
        .ARST_N                    ( LANECTRL_ADDR_CMD_0_ARST_N ),
        .RX_SYNC_RST               ( LANECTRL_ADDR_CMD_0_RX_SYNC_RST ),
        .TX_SYNC_RST               ( LANECTRL_ADDR_CMD_0_TX_SYNC_RST ),
        .HS_IO_CLK                 ( HS_IO_CLK ),
        .TX_DQS_270                ( LANECTRL_ADDR_CMD_0_TX_DQS_270 ),
        .TX_DATA_0                 ( TX_DATA_0_net_4 ),
        .TX_DATA_1                 ( TX_DATA_1_net_1 ),
        .OE_DATA_0                 ( OE_DATA_0_const_net_3 ),
        .OE_DATA_1                 ( OE_DATA_1_const_net_1 ),
        .DELAY_LINE_MOVE_0         ( IOD_TRAINING_0_CMD_DELAY_LINE_MOVE ),
        .DELAY_LINE_MOVE_1         ( IOD_TRAINING_0_CMD_DELAY_LINE_MOVE ),
        .DELAY_LINE_DIRECTION_0    ( IOD_TRAINING_0_CMD_DELAY_LINE_DIRECTION ),
        .DELAY_LINE_DIRECTION_1    ( IOD_TRAINING_0_CMD_DELAY_LINE_DIRECTION ),
        .DELAY_LINE_LOAD_0         ( IOD_TRAINING_0_CMD_DELAY_LINE_LOAD ),
        .DELAY_LINE_LOAD_1         ( IOD_TRAINING_0_CMD_DELAY_LINE_LOAD ),
        .FAB_CLK                   ( SYS_CLK ),
        .ODT_EN_0                  ( GND_net ), // tied to 1'b0 from definition
        .ODT_EN_1                  ( GND_net ), // tied to 1'b0 from definition
        // Outputs
        .DELAY_LINE_OUT_OF_RANGE_0 (  ),
        .DELAY_LINE_OUT_OF_RANGE_1 (  ),
        .PAD_O                     ( BA_net_0 ) 
        );

//--------PF_DDR4_SS_DDRPHY_BLK_IOD_BCLK_TRAINING_PF_IOD   -   Actel:SgCore:PF_IOD:1.0.218
PF_DDR4_SS_DDRPHY_BLK_IOD_BCLK_TRAINING_PF_IOD IOD_BCLK_TRAINING(
        // Inputs
        .ARST_N                    ( VCC_net ), // tied to 1'b1 from definition
        .RX_SYNC_RST               ( VCC_net ), // tied to 1'b1 from definition
        .TX_SYNC_RST               ( VCC_net ), // tied to 1'b1 from definition
        .HS_IO_CLK                 ( HS_IO_CLK ),
        .EYE_MONITOR_CLEAR_FLAGS_0 ( IOD_TRAINING_0_BCLK_EYE_MONITOR_CLR_FLAGS ),
        .DELAY_LINE_MOVE_0         ( GND_net ),
        .DELAY_LINE_DIRECTION_0    ( GND_net ),
        .DELAY_LINE_LOAD_0         ( GND_net ),
        .FAB_CLK                   ( SYS_CLK ),
        .ODT_EN_0                  ( GND_net ), // tied to 1'b0 from definition
        // Outputs
        .DELAY_LINE_OUT_OF_RANGE_0 (  ),
        .EYE_MONITOR_EARLY_0       ( IOD_BCLK_TRAINING_EYE_MONITOR_EARLY_0 ),
        .EYE_MONITOR_LATE_0        ( IOD_BCLK_TRAINING_EYE_MONITOR_LATE_0 ),
        .RX_DATA_0                 ( RX_DATA_0_net_1 ) 
        );

//--------PF_DDR4_SS_DDRPHY_BLK_IOD_BG_PF_IOD   -   Actel:SgCore:PF_IOD:1.0.218
PF_DDR4_SS_DDRPHY_BLK_IOD_BG_PF_IOD IOD_BG(
        // Inputs
        .ARST_N                    ( LANECTRL_ADDR_CMD_0_ARST_N ),
        .RX_SYNC_RST               ( LANECTRL_ADDR_CMD_0_RX_SYNC_RST ),
        .TX_SYNC_RST               ( LANECTRL_ADDR_CMD_0_TX_SYNC_RST ),
        .HS_IO_CLK                 ( HS_IO_CLK ),
        .TX_DQS_270                ( LANECTRL_ADDR_CMD_0_TX_DQS_270 ),
        .TX_DATA_0                 ( TX_DATA_0_net_5 ),
        .TX_DATA_1                 ( TX_DATA_1_net_2 ),
        .OE_DATA_0                 ( OE_DATA_0_const_net_4 ),
        .OE_DATA_1                 ( OE_DATA_1_const_net_2 ),
        .DELAY_LINE_MOVE_0         ( IOD_TRAINING_0_CMD_DELAY_LINE_MOVE ),
        .DELAY_LINE_MOVE_1         ( IOD_TRAINING_0_CMD_DELAY_LINE_MOVE ),
        .DELAY_LINE_DIRECTION_0    ( IOD_TRAINING_0_CMD_DELAY_LINE_DIRECTION ),
        .DELAY_LINE_DIRECTION_1    ( IOD_TRAINING_0_CMD_DELAY_LINE_DIRECTION ),
        .DELAY_LINE_LOAD_0         ( IOD_TRAINING_0_CMD_DELAY_LINE_LOAD ),
        .DELAY_LINE_LOAD_1         ( IOD_TRAINING_0_CMD_DELAY_LINE_LOAD ),
        .FAB_CLK                   ( SYS_CLK ),
        .ODT_EN_0                  ( GND_net ), // tied to 1'b0 from definition
        .ODT_EN_1                  ( GND_net ), // tied to 1'b0 from definition
        // Outputs
        .DELAY_LINE_OUT_OF_RANGE_0 (  ),
        .DELAY_LINE_OUT_OF_RANGE_1 (  ),
        .PAD_O                     ( BG_net_0 ) 
        );

//--------PF_DDR4_SS_DDRPHY_BLK_IOD_CAS_N_PF_IOD   -   Actel:SgCore:PF_IOD:1.0.218
PF_DDR4_SS_DDRPHY_BLK_IOD_CAS_N_PF_IOD IOD_CAS_N(
        // Inputs
        .ARST_N                    ( LANECTRL_ADDR_CMD_0_ARST_N ),
        .RX_SYNC_RST               ( LANECTRL_ADDR_CMD_0_RX_SYNC_RST ),
        .TX_SYNC_RST               ( LANECTRL_ADDR_CMD_0_TX_SYNC_RST ),
        .HS_IO_CLK                 ( HS_IO_CLK ),
        .TX_DQS_270                ( LANECTRL_ADDR_CMD_0_TX_DQS_270 ),
        .TX_DATA_0                 ( TX_DATA_0_net_6 ),
        .OE_DATA_0                 ( OE_DATA_0_const_net_5 ),
        .DELAY_LINE_MOVE_0         ( IOD_TRAINING_0_CMD_DELAY_LINE_MOVE ),
        .DELAY_LINE_DIRECTION_0    ( IOD_TRAINING_0_CMD_DELAY_LINE_DIRECTION ),
        .DELAY_LINE_LOAD_0         ( IOD_TRAINING_0_CMD_DELAY_LINE_LOAD ),
        .FAB_CLK                   ( SYS_CLK ),
        .ODT_EN_0                  ( GND_net ), // tied to 1'b0 from definition
        // Outputs
        .DELAY_LINE_OUT_OF_RANGE_0 (  ),
        .PAD_O                     ( CAS_N_net_0 ) 
        );

//--------PF_DDR4_SS_DDRPHY_BLK_IOD_CKE_PF_IOD   -   Actel:SgCore:PF_IOD:1.0.218
PF_DDR4_SS_DDRPHY_BLK_IOD_CKE_PF_IOD IOD_CKE(
        // Inputs
        .ARST_N                    ( LANECTRL_ADDR_CMD_0_ARST_N ),
        .RX_SYNC_RST               ( LANECTRL_ADDR_CMD_0_RX_SYNC_RST ),
        .TX_SYNC_RST               ( LANECTRL_ADDR_CMD_0_TX_SYNC_RST ),
        .HS_IO_CLK                 ( HS_IO_CLK ),
        .TX_DQS_270                ( LANECTRL_ADDR_CMD_0_TX_DQS_270 ),
        .TX_DATA_0                 ( TX_DATA_0_net_7 ),
        .OE_DATA_0                 ( OE_DATA_0_const_net_6 ),
        .DELAY_LINE_MOVE_0         ( GND_net ),
        .DELAY_LINE_DIRECTION_0    ( GND_net ),
        .DELAY_LINE_LOAD_0         ( GND_net ),
        .FAB_CLK                   ( SYS_CLK ),
        .ODT_EN_0                  ( GND_net ), // tied to 1'b0 from definition
        // Outputs
        .DELAY_LINE_OUT_OF_RANGE_0 (  ),
        .PAD_O                     ( CKE_net_0 ) 
        );

//--------PF_DDR4_SS_DDRPHY_BLK_IOD_CS_N_PF_IOD   -   Actel:SgCore:PF_IOD:1.0.218
PF_DDR4_SS_DDRPHY_BLK_IOD_CS_N_PF_IOD IOD_CS_N(
        // Inputs
        .ARST_N                    ( LANECTRL_ADDR_CMD_0_ARST_N ),
        .RX_SYNC_RST               ( LANECTRL_ADDR_CMD_0_RX_SYNC_RST ),
        .TX_SYNC_RST               ( LANECTRL_ADDR_CMD_0_TX_SYNC_RST ),
        .HS_IO_CLK                 ( HS_IO_CLK ),
        .TX_DQS_270                ( LANECTRL_ADDR_CMD_0_TX_DQS_270 ),
        .TX_DATA_0                 ( TX_DATA_0_net_8 ),
        .OE_DATA_0                 ( OE_DATA_0_const_net_7 ),
        .DELAY_LINE_MOVE_0         ( IOD_TRAINING_0_CMD_DELAY_LINE_MOVE ),
        .DELAY_LINE_DIRECTION_0    ( IOD_TRAINING_0_CMD_DELAY_LINE_DIRECTION ),
        .DELAY_LINE_LOAD_0         ( IOD_TRAINING_0_CMD_DELAY_LINE_LOAD ),
        .FAB_CLK                   ( SYS_CLK ),
        .ODT_EN_0                  ( GND_net ), // tied to 1'b0 from definition
        // Outputs
        .DELAY_LINE_OUT_OF_RANGE_0 (  ),
        .PAD_O                     ( CS_N_net_0 ) 
        );

//--------PF_DDR4_SS_DDRPHY_BLK_IOD_ODT_PF_IOD   -   Actel:SgCore:PF_IOD:1.0.218
PF_DDR4_SS_DDRPHY_BLK_IOD_ODT_PF_IOD IOD_ODT(
        // Inputs
        .ARST_N                    ( LANECTRL_ADDR_CMD_0_ARST_N ),
        .RX_SYNC_RST               ( LANECTRL_ADDR_CMD_0_RX_SYNC_RST ),
        .TX_SYNC_RST               ( LANECTRL_ADDR_CMD_0_TX_SYNC_RST ),
        .HS_IO_CLK                 ( HS_IO_CLK ),
        .TX_DQS_270                ( LANECTRL_ADDR_CMD_0_TX_DQS_270 ),
        .TX_DATA_0                 ( TX_DATA_0_net_9 ),
        .OE_DATA_0                 ( OE_DATA_0_const_net_8 ),
        .DELAY_LINE_MOVE_0         ( IOD_TRAINING_0_CMD_DELAY_LINE_MOVE ),
        .DELAY_LINE_DIRECTION_0    ( IOD_TRAINING_0_CMD_DELAY_LINE_DIRECTION ),
        .DELAY_LINE_LOAD_0         ( IOD_TRAINING_0_CMD_DELAY_LINE_LOAD ),
        .FAB_CLK                   ( SYS_CLK ),
        .ODT_EN_0                  ( GND_net ), // tied to 1'b0 from definition
        // Outputs
        .DELAY_LINE_OUT_OF_RANGE_0 (  ),
        .PAD_O                     ( ODT_net_0 ) 
        );

//--------PF_DDR4_SS_DDRPHY_BLK_IOD_RAS_N_PF_IOD   -   Actel:SgCore:PF_IOD:1.0.218
PF_DDR4_SS_DDRPHY_BLK_IOD_RAS_N_PF_IOD IOD_RAS_N(
        // Inputs
        .ARST_N                    ( LANECTRL_ADDR_CMD_0_ARST_N ),
        .RX_SYNC_RST               ( LANECTRL_ADDR_CMD_0_RX_SYNC_RST ),
        .TX_SYNC_RST               ( LANECTRL_ADDR_CMD_0_TX_SYNC_RST ),
        .HS_IO_CLK                 ( HS_IO_CLK ),
        .TX_DQS_270                ( LANECTRL_ADDR_CMD_0_TX_DQS_270 ),
        .TX_DATA_0                 ( TX_DATA_0_net_10 ),
        .OE_DATA_0                 ( OE_DATA_0_const_net_9 ),
        .DELAY_LINE_MOVE_0         ( IOD_TRAINING_0_CMD_DELAY_LINE_MOVE ),
        .DELAY_LINE_DIRECTION_0    ( IOD_TRAINING_0_CMD_DELAY_LINE_DIRECTION ),
        .DELAY_LINE_LOAD_0         ( IOD_TRAINING_0_CMD_DELAY_LINE_LOAD ),
        .FAB_CLK                   ( SYS_CLK ),
        .ODT_EN_0                  ( GND_net ), // tied to 1'b0 from definition
        // Outputs
        .DELAY_LINE_OUT_OF_RANGE_0 (  ),
        .PAD_O                     ( RAS_N_net_0 ) 
        );

//--------PF_DDR4_SS_DDRPHY_BLK_IOD_REF_CLK_TRAINING_PF_IOD   -   Actel:SgCore:PF_IOD:1.0.218
PF_DDR4_SS_DDRPHY_BLK_IOD_REF_CLK_TRAINING_PF_IOD IOD_REF_CLK_TRAINING(
        // Inputs
        .RX_P_0                    ( OB_DIFF_CK0_Y ),
        .HS_IO_CLK                 ( HS_IO_CLK ),
        .EYE_MONITOR_CLEAR_FLAGS_0 ( IOD_TRAINING_0_REFCLK_EYE_MONITOR_CLR_FLAGS ),
        .DELAY_LINE_MOVE_0         ( IOD_TRAINING_0_REFCLK_DELAY_LINE_MOVE ),
        .DELAY_LINE_DIRECTION_0    ( IOD_TRAINING_0_REFCLK_DELAY_LINE_DIRECTION ),
        .DELAY_LINE_LOAD_0         ( IOD_TRAINING_0_REFCLK_DELAY_LINE_LOAD ),
        .FAB_CLK                   ( SYS_CLK ),
        .ODT_EN_0                  ( GND_net ), // tied to 1'b0 from definition
        // Outputs
        .DELAY_LINE_OUT_OF_RANGE_0 (  ),
        .EYE_MONITOR_EARLY_0       ( IOD_REF_CLK_TRAINING_EYE_MONITOR_EARLY_0 ),
        .EYE_MONITOR_LATE_0        ( IOD_REF_CLK_TRAINING_EYE_MONITOR_LATE_0 ),
        .RX_DATA_0                 ( RX_DATA_0_net_2 ) 
        );

//--------PF_DDR4_SS_DDRPHY_BLK_IOD_RESET_N_PF_IOD   -   Actel:SgCore:PF_IOD:1.0.218
PF_DDR4_SS_DDRPHY_BLK_IOD_RESET_N_PF_IOD IOD_RESET_N(
        // Inputs
        .ARST_N                    ( LANECTRL_ADDR_CMD_0_ARST_N ),
        .RX_SYNC_RST               ( LANECTRL_ADDR_CMD_0_RX_SYNC_RST ),
        .TX_SYNC_RST               ( LANECTRL_ADDR_CMD_0_TX_SYNC_RST ),
        .HS_IO_CLK                 ( HS_IO_CLK ),
        .TX_DQS_270                ( LANECTRL_ADDR_CMD_0_TX_DQS_270 ),
        .TX_DATA_0                 ( TX_DATA_0_net_11 ),
        .OE_DATA_0                 ( OE_DATA_0_const_net_10 ),
        .DELAY_LINE_MOVE_0         ( GND_net ),
        .DELAY_LINE_DIRECTION_0    ( GND_net ),
        .DELAY_LINE_LOAD_0         ( GND_net ),
        .FAB_CLK                   ( SYS_CLK ),
        .ODT_EN_0                  ( GND_net ), // tied to 1'b0 from definition
        // Outputs
        .DELAY_LINE_OUT_OF_RANGE_0 (  ),
        .PAD_O                     ( RESET_N_net_0 ) 
        );

//--------COREDDR_TIP   -   Actel:DirectCore:COREDDR_TIP:2.1.101
COREDDR_TIP #( 
        .FAMILY             ( 26 ),
        .FIFO_ADDRESS_WIDTH ( 7 ),
        .FIFO_DEPTH         ( 2 ),
        .IOG_DQ_WIDTH_L0    ( 8 ),
        .IOG_DQ_WIDTH_L1    ( 8 ),
        .IOG_DQ_WIDTH_L2    ( 8 ),
        .IOG_DQ_WIDTH_L3    ( 8 ),
        .IOG_DQ_WIDTH_L4    ( 8 ),
        .IOG_DQ_WIDTH_L5    ( 8 ),
        .IOG_DQ_WIDTH_L6    ( 8 ),
        .IOG_DQ_WIDTH_L7    ( 8 ),
        .IOG_DQ_WIDTH_L8    ( 8 ),
        .IOG_DQS_LANES      ( 4 ),
        .NUM_BCLKS          ( 1 ),
        .PIPELINE           ( 1 ),
        .SIM_TRAINING       ( 0 ) )
IOD_TRAINING_0(
        // Inputs
        .SCLK                          ( SYS_CLK ),
        .RESET_N                       ( SYS_RST_N ),
        .DFI_INIT_START                ( DFI_INIT_START ),
        .DFI_RDLVL_CS_0_N              ( DFI_RDLVL_CS_N ),
        .DFI_RDLVL_CS_1_N              ( VCC_net ),
        .DFI_WRLVL_CS_0_N              ( DFI_WRLVL_CS_N ),
        .DFI_WRLVL_CS_1_N              ( VCC_net ),
        .DFI_RDDATA_CS_0_N_P0          ( DFI_RDDATA_CS_N_P0 ),
        .DFI_RDDATA_CS_0_N_P1          ( DFI_RDDATA_CS_N_P1 ),
        .DFI_RDDATA_CS_0_N_P2          ( DFI_RDDATA_CS_N_P2 ),
        .DFI_RDDATA_CS_0_N_P3          ( DFI_RDDATA_CS_N_P3 ),
        .DFI_RDDATA_CS_1_N_P0          ( GND_net ),
        .DFI_RDDATA_CS_1_N_P1          ( GND_net ),
        .DFI_RDDATA_CS_1_N_P2          ( GND_net ),
        .DFI_RDDATA_CS_1_N_P3          ( GND_net ),
        .DFI_WRDATA_CS_0_N_P0          ( DFI_WRDATA_CS_N_P0 ),
        .DFI_WRDATA_CS_0_N_P1          ( DFI_WRDATA_CS_N_P1 ),
        .DFI_WRDATA_CS_0_N_P2          ( DFI_WRDATA_CS_N_P2 ),
        .DFI_WRDATA_CS_0_N_P3          ( DFI_WRDATA_CS_N_P3 ),
        .DFI_WRDATA_CS_1_N_P0          ( GND_net ),
        .DFI_WRDATA_CS_1_N_P1          ( GND_net ),
        .DFI_WRDATA_CS_1_N_P2          ( GND_net ),
        .DFI_WRDATA_CS_1_N_P3          ( GND_net ),
        .DFI_RDLVL_EN                  ( DFI_RDLVL_EN ),
        .DFI_RDLVL_GATE_EN             ( DFI_RDLVL_GATE_EN ),
        .DFI_WRDATA_EN_P0              ( DFI_WRDATA_EN_P0_slice_0 ),
        .DFI_WRDATA_EN_P1              ( DFI_WRDATA_EN_P1_slice_0 ),
        .DFI_WRDATA_EN_P2              ( DFI_WRDATA_EN_P2_slice_0 ),
        .DFI_WRDATA_EN_P3              ( DFI_WRDATA_EN_P3_slice_0 ),
        .DFI_WRLVL_EN                  ( DFI_WRLVL_EN ),
        .DFI_WRLVL_STROBE              ( DFI_WRLVL_STROBE ),
        .BCLK_EYE_MONITOR_EARLY        ( IOD_BCLK_TRAINING_EYE_MONITOR_EARLY_0 ),
        .BCLK_EYE_MONITOR_LATE         ( IOD_BCLK_TRAINING_EYE_MONITOR_LATE_0 ),
        .BURST_DETECT                  ( BURST_DETECT_net_0 ),
        .REFCLK_EYE_MONITOR_EARLY      ( IOD_REF_CLK_TRAINING_EYE_MONITOR_EARLY_0 ),
        .REFCLK_EYE_MONITOR_LATE       ( IOD_REF_CLK_TRAINING_EYE_MONITOR_LATE_0 ),
        .RX_OUT_OF_RANGE               ( RX_OUT_OF_RANGE_net_0 ),
        .TWO_RANKS                     ( GND_net ),
        .TX_OUT_OF_RANGE               ( TX_OUT_OF_RANGE_net_0 ),
        .PADDR                         ( PADDR ),
        .PENABLE                       ( PENABLE ),
        .PSEL                          ( PSEL ),
        .PWDATA                        ( PWDATA ),
        .PWRITE                        ( PWRITE ),
        .TRAINING_PATTERN              ( TRAINING_PATTERN_const_net_0 ),
        .DLL_DLY_DIFF                  ( DLL_DLY_DIFF ),
        .VREF_OUT_OF_RANGE             (  ),
        .DFI_CTRLUPD_REQ               ( DFI_CTRLUPD_REQ ),
        .DFI_RDDATA_EN_P0              ( DFI_RDDATA_EN_P0_slice_0 ),
        .DFI_RDDATA_EN_P1              ( DFI_RDDATA_EN_P1_slice_0 ),
        .DFI_RDDATA_EN_P2              ( DFI_RDDATA_EN_P2_slice_0 ),
        .DFI_RDDATA_EN_P3              ( DFI_RDDATA_EN_P3_slice_0 ),
        .IOG_RDDATA                    ( IOG_RDDATA_net_0 ),
        .IOG_RDDATA_VALID              ( IOG_RDDATA_VALID_net_0 ),
        .PAD_RDDATA                    ( PAD_RDDATA_net_0 ),
        .DQSW_EYE_MONITOR_EARLY        ( DQSW_EYE_MONITOR_EARLY_net_0 ),
        .DQSW_EYE_MONITOR_LATE         ( DQSW_EYE_MONITOR_LATE_net_0 ),
        .DQSW270_EYE_MONITOR_EARLY     ( DQSW270_EYE_MONITOR_EARLY_net_0 ),
        .DQSW270_EYE_MONITOR_LATE      ( DQSW270_EYE_MONITOR_LATE_net_0 ),
        .CMD_EYE_MONITOR_EARLY         ( IOD_A_12_EYE_MONITOR_EARLY_0 ),
        .CMD_EYE_MONITOR_LATE          ( IOD_A_12_EYE_MONITOR_LATE_0 ),
        .REFCLK_IGEAR_RX8              ( IOD_REF_CLK_TRAINING_RX_DATA_06to6 ),
        .DQSW270_IGEAR_RX8             ( DQSW270_IGEAR_RX8_net_0 ),
        .DQSW_DELAY_LINE_OOR           ( DQSW_DELAY_LINE_OOR_net_0 ),
        .DQSW270_DELAY_LINE_OOR        ( DQSW270_DELAY_LINE_OOR_net_0 ),
        .PLL_LOCK                      ( PLL_LOCK ),
        .DFI_WRDATA_MASK_P0            (  ),
        .DFI_WRDATA_MASK_P1            (  ),
        .DFI_WRDATA_MASK_P2            (  ),
        .DFI_WRDATA_MASK_P3            (  ),
        .DFI_ADDRESS_P0                ( DFI_ADDRESS_P0_net_0 ),
        .DFI_ADDRESS_P1                ( DFI_ADDRESS_P1_net_0 ),
        .DFI_ADDRESS_P2                ( DFI_ADDRESS_P2_net_0 ),
        .DFI_ADDRESS_P3                ( DFI_ADDRESS_P3_net_0 ),
        .BCLK_IGEAR_RX                 ( BCLK_IGEAR_RX_net_0 ),
        .CMD_IGEAR_RX8                 ( IOD_A_12_RX_DATA_03to3 ),
        .DQSW270_IGEAR_RX              ( DQSW270_IGEAR_RX_net_0 ),
        .DQSW_IGEAR_RX                 ( DQSW_IGEAR_RX_net_0 ),
        .SKIP_DQSW_TRN                 ( SKIP_DQSW_TRN ),
        .SKIP_BCLK_TRN                 ( SKIP_BCLK_TRN ),
        .SKIP_CA_TRN                   ( SKIP_CA_TRN ),
        .SKIP_WRLVL_TRN                ( SKIP_WRLVL_TRN ),
        .SKIP_RDLVL_TRN                ( SKIP_RDLVL_TRN ),
        .BCLK_VCOPHS_OFFSET            ( BCLK_VCOPHS_OFFSET ),
        .ADDR_VCOPHS_OFFSET            ( ADDR_VCOPHS_OFFSET ),
        .WRLVL_TAP_OFFSET              ( WRLVL_TAP_OFFSET ),
        .CAL_INIT_ACK                  ( CAL_INIT_ACK ),
        .SKIP_VREF_TRAINING            ( SKIP_VREF_TRAINING ),
        .PCLK                          ( PCLK ),
        .VREF_MR6_VALUE                ( VREF_MR6_VALUE ),
        .CTRLR_READY_IN                ( CTRLR_READY_IN ),
        .IOG_DQ_TXDATA_IN              ( IOG_DQ_TXDATA_IN_net_0 ),
        .IOG_DM_TXDATA_IN              ( IOG_DM_TXDATA_IN_net_0 ),
        .CAL_L_BUSY                    ( CAL_L_BUSY ),
        .CAL_L_D_REQ                   ( CAL_L_D_REQ ),
        .CAL_L_DATAOUT                 ( CAL_L_DATAOUT ),
        .CAL_L_R_VALID                 ( CAL_L_R_VALID ),
        .ADDR_WAIT_COUNT               ( ADDR_WAIT_COUNT ),
        .WRCAL_WRITE_COUNTER_VALUE     ( WRCAL_WRITE_COUNTER_VALUE ),
        .RDGATE_MIN_READS_THRESHOLD    ( RDGATE_MIN_READS_THRESHOLD ),
        .DFI_RESET_N_P0                ( DFI_RESET_N_P0 ),
        .DFI_RESET_N_P1                ( DFI_RESET_N_P1 ),
        .DFI_RESET_N_P2                ( DFI_RESET_N_P2 ),
        .DFI_RESET_N_P3                ( DFI_RESET_N_P3 ),
        .DFI_BANK_P0                   ( DFI_BANK_P0_net_0 ),
        .DFI_BANK_P1                   ( DFI_BANK_P1_net_0 ),
        .DFI_BANK_P2                   ( DFI_BANK_P2_net_0 ),
        .DFI_BANK_P3                   ( DFI_BANK_P3_net_0 ),
        .DFI_CS_N_P0                   ( DFI_CS_N_P0 ),
        .DFI_CS_N_P1                   ( DFI_CS_N_P1 ),
        .DFI_CS_N_P2                   ( DFI_CS_N_P2 ),
        .DFI_CS_N_P3                   ( DFI_CS_N_P3 ),
        .DFI_ODT_P0                    ( DFI_ODT_P0 ),
        .DFI_ODT_P1                    ( DFI_ODT_P1 ),
        .DFI_ODT_P2                    ( DFI_ODT_P2 ),
        .DFI_ODT_P3                    ( DFI_ODT_P3 ),
        .DFI_CKE_P0                    ( DFI_CKE_P0 ),
        .DFI_CKE_P1                    ( DFI_CKE_P1 ),
        .DFI_CKE_P2                    ( DFI_CKE_P2 ),
        .DFI_CKE_P3                    ( DFI_CKE_P3 ),
        .DFI_RAS_N_P0                  ( DFI_RAS_N_P0 ),
        .DFI_RAS_N_P1                  ( DFI_RAS_N_P1 ),
        .DFI_RAS_N_P2                  ( DFI_RAS_N_P2 ),
        .DFI_RAS_N_P3                  ( DFI_RAS_N_P3 ),
        .DFI_CAS_N_P0                  ( DFI_CAS_N_P0 ),
        .DFI_CAS_N_P1                  ( DFI_CAS_N_P1 ),
        .DFI_CAS_N_P2                  ( DFI_CAS_N_P2 ),
        .DFI_CAS_N_P3                  ( DFI_CAS_N_P3 ),
        .DFI_WE_N_P0                   ( DFI_WE_N_P0 ),
        .DFI_WE_N_P1                   ( DFI_WE_N_P1 ),
        .DFI_WE_N_P2                   ( DFI_WE_N_P2 ),
        .DFI_WE_N_P3                   ( DFI_WE_N_P3 ),
        .DFI_ACT_N_P0                  ( DFI_ACT_N_P0 ),
        .DFI_ACT_N_P1                  ( DFI_ACT_N_P1 ),
        .DFI_ACT_N_P2                  ( DFI_ACT_N_P2 ),
        .DFI_ACT_N_P3                  ( DFI_ACT_N_P3 ),
        .DFI_BG_P0                     ( DFI_BG_P0_net_0 ),
        .DFI_BG_P1                     ( DFI_BG_P1_net_0 ),
        .DFI_BG_P2                     ( DFI_BG_P2_net_0 ),
        .DFI_BG_P3                     ( DFI_BG_P3_net_0 ),
        // Outputs
        .DFI_INIT_COMPLETE             ( DFI_INIT_COMPLETE_net_0 ),
        .DFI_RDLVL_RESP                ( DFI_RDLVL_RESP_net_0 ),
        .DFI_TRAINING_COMPLETE         ( DFI_TRAINING_COMPLETE_net_0 ),
        .DFI_WRLVL_RESP                ( DFI_WRLVL_RESP_net_0 ),
        .BCLK_EYE_MONITOR_CLR_FLAGS    ( IOD_TRAINING_0_BCLK_EYE_MONITOR_CLR_FLAGS ),
        .CLK_SEL                       ( CLK_SEL_net_0 ),
        .DELAY_LINE_SEL_RD             ( DELAY_LINE_SEL_RD_net_0 ),
        .DIRECTION                     ( DIRECTION_net_0 ),
        .IOG_OE_P0                     ( IOG_OE_P0_net_0 ),
        .IOG_OE_P1                     ( IOG_OE_P1_net_0 ),
        .IOG_OE_P2                     ( IOG_OE_P2_net_0 ),
        .IOG_OE_P3                     ( IOG_OE_P3_net_0 ),
        .DQS_OE_P0                     ( DQS_OE_P0_net_0 ),
        .DQS_OE_P1                     ( DQS_OE_P1_net_0 ),
        .DQS_OE_P2                     ( DQS_OE_P2_net_0 ),
        .DQS_OE_P3                     ( DQS_OE_P3_net_0 ),
        .DM_OE_P0                      ( DM_OE_P0_net_0 ),
        .DM_OE_P1                      ( DM_OE_P1_net_0 ),
        .DM_OE_P2                      ( DM_OE_P2_net_0 ),
        .DM_OE_P3                      ( DM_OE_P3_net_0 ),
        .LOAD                          ( LOAD_net_0 ),
        .MOVE                          ( MOVE_net_0 ),
        .REFCLK_EYE_MONITOR_CLR_FLAGS  ( IOD_TRAINING_0_REFCLK_EYE_MONITOR_CLR_FLAGS ),
        .PRDATA                        ( APB_DEBUG_PRDATA ),
        .PREADY                        ( APB_DEBUG_PREADY ),
        .ODT_DYN_LANE                  ( ODT_DYN_LANE_net_0 ),
        .CODE_UPDATE                   ( CODE_UPDATE_net_0 ),
        .LOADPHS_B                     ( LOADPHS_B_net_0 ),
        .VCO_PHSEL_BCLK_SEL            ( VCO_PHSEL_BCLK_SEL_net_0 ),
        .VCO_PHSEL_REFCLK_SEL          ( VCO_PHSEL_REFCLK_SEL_net_0 ),
        .VCO_PHSEL_ROTATE              ( VCO_PHSEL_ROTATE_net_0 ),
        .VREF_DIRECTION                (  ),
        .VREF_MOVE                     (  ),
        .VREF_RELOAD                   (  ),
        .DFI_RDDATA_W0                 ( DFI_RDDATA_W0_net_0 ),
        .DFI_RDDATA_W1                 ( DFI_RDDATA_W1_net_0 ),
        .DFI_RDDATA_W2                 ( DFI_RDDATA_W2_net_0 ),
        .DFI_RDDATA_W3                 ( DFI_RDDATA_W3_net_0 ),
        .DFI_RDDATA_VALID_W0           ( DFI_RDDATA_VALID_W0_net_0 ),
        .DFI_RDDATA_VALID_W1           ( DFI_RDDATA_VALID_W1_net_0 ),
        .DFI_RDDATA_VALID_W2           ( DFI_RDDATA_VALID_W2_net_0 ),
        .DFI_RDDATA_VALID_W3           ( DFI_RDDATA_VALID_W3_net_0 ),
        .IOG_RDDATA_EN_P0_P            ( IOG_RDDATA_EN_P0_P_net_0 ),
        .IOG_RDDATA_EN_P0_N            ( IOG_RDDATA_EN_P0_N_net_0 ),
        .IOG_RDDATA_EN_P1_P            ( IOG_RDDATA_EN_P1_P_net_0 ),
        .IOG_RDDATA_EN_P1_N            ( IOG_RDDATA_EN_P1_N_net_0 ),
        .IOG_RDDATA_EN_P2_P            ( IOG_RDDATA_EN_P2_P_net_0 ),
        .IOG_RDDATA_EN_P2_N            ( IOG_RDDATA_EN_P2_N_net_0 ),
        .IOG_RDDATA_EN_P3_P            ( IOG_RDDATA_EN_P3_P_net_0 ),
        .IOG_RDDATA_EN_P3_N            ( IOG_RDDATA_EN_P3_N_net_0 ),
        .RD_TRAINING_ERROR             (  ),
        .DQSW_EYE_MONITOR_CLR_FLAGS    ( DQSW_EYE_MONITOR_CLR_FLAGS_net_0 ),
        .DQSW270_EYE_MONITOR_CLR_FLAGS ( DQSW270_EYE_MONITOR_CLR_FLAGS_net_0 ),
        .DQSW_DELAY_LINE_LOAD          ( DQSW_DELAY_LINE_LOAD_net_0 ),
        .DQSW_DELAY_LINE_MOVE          ( DQSW_DELAY_LINE_MOVE_net_0 ),
        .DQSW_DELAY_LINE_DIRECTION     ( DQSW_DELAY_LINE_DIRECTION_net_0 ),
        .DQSW270_DELAY_LINE_LOAD       ( DQSW270_DELAY_LINE_LOAD_net_0 ),
        .DQSW270_DELAY_LINE_MOVE       ( DQSW270_DELAY_LINE_MOVE_net_0 ),
        .DQSW270_DELAY_LINE_DIRECTION  ( DQSW270_DELAY_LINE_DIRECTION_net_0 ),
        .REFCLK_DELAY_LINE_LOAD        ( IOD_TRAINING_0_REFCLK_DELAY_LINE_LOAD ),
        .REFCLK_DELAY_LINE_MOVE        ( IOD_TRAINING_0_REFCLK_DELAY_LINE_MOVE ),
        .REFCLK_DELAY_LINE_DIRECTION   ( IOD_TRAINING_0_REFCLK_DELAY_LINE_DIRECTION ),
        .CMD_EYE_MONITOR_CLR_FLAGS     ( IOD_TRAINING_0_CMD_EYE_MONITOR_CLR_FLAGS ),
        .CMD_DELAY_LINE_LOAD           ( IOD_TRAINING_0_CMD_DELAY_LINE_LOAD ),
        .CMD_DELAY_LINE_MOVE           ( IOD_TRAINING_0_CMD_DELAY_LINE_MOVE ),
        .CMD_DELAY_LINE_DIRECTION      ( IOD_TRAINING_0_CMD_DELAY_LINE_DIRECTION ),
        .VCO_PHSEL_BCLK90_SEL          ( VCO_PHSEL_BCLK90_SEL_net_0 ),
        .DQSW_SELA                     ( DQSW_SELA_net_0 ),
        .CMD_OE                        ( IOD_TRAINING_0_CMD_OE ),
        .CMD_DELAY_LINE_MOVE_TRN       ( IOD_TRAINING_0_CMD_DELAY_LINE_MOVE_TRN ),
        .INIT_PAUSE                    ( INIT_PAUSE_net_0 ),
        .INIT_RESET                    ( SYNC_SYS_RST_N_net_0 ),
        .IOG_WRDATA_MASK_P0            ( IOG_WRDATA_MASK_P0_net_0 ),
        .IOG_WRDATA_MASK_P1            ( IOG_WRDATA_MASK_P1_net_0 ),
        .IOG_WRDATA_MASK_P2            ( IOG_WRDATA_MASK_P2_net_0 ),
        .IOG_WRDATA_MASK_P3            ( IOG_WRDATA_MASK_P3_net_0 ),
        .IOG_ADDRESS_P0                ( IOG_ADDRESS_P0_net_0 ),
        .IOG_ADDRESS_P1                ( IOG_ADDRESS_P1_net_0 ),
        .IOG_ADDRESS_P2                ( IOG_ADDRESS_P2_net_0 ),
        .IOG_ADDRESS_P3                ( IOG_ADDRESS_P3_net_0 ),
        .CMD_RESET_LANE                ( IOD_TRAINING_0_CMD_RESET_LANE ),
        .CAL_INIT_MR_W_REQ             ( CAL_INIT_MR_W_REQ_net_0 ),
        .CAL_INIT_MR_ADDR              ( CAL_INIT_MR_ADDR_net_0 ),
        .CAL_INIT_MR_WR_DATA           ( CAL_INIT_MR_WR_DATA_net_0 ),
        .CAL_INIT_MR_WR_MASK           ( CAL_INIT_MR_WR_MASK_net_0 ),
        .CAL_INIT_CS                   ( CAL_INIT_CS_net_0 ),
        .CTRLR_READY_OUT               ( CTRLR_READY_OUT_net_0 ),
        .IOG_DQ_TXDATA_OUT             ( IOG_DQ_TXDATA_OUT_net_0 ),
        .IOG_DM_TXDATA_OUT             ( IOG_DM_TXDATA_OUT_net_0 ),
        .CAL_L_R_REQ                   ( CAL_L_R_REQ_net_0 ),
        .CAL_L_W_REQ                   ( CAL_L_W_REQ_net_0 ),
        .CAL_L_DATAIN                  ( CAL_L_DATAIN_net_0 ),
        .CAL_L_DM_IN                   ( CAL_L_DM_IN_net_0 ),
        .CAL_SELECT                    ( CAL_SELECT_net_0 ),
        .ITER_COUNT                    ( ITER_COUNT_net_0 ),
        .DFI_RESET_N_P0_OUT            ( IOD_TRAINING_0_DFI_RESET_N_P0_OUT ),
        .DFI_RESET_N_P1_OUT            ( IOD_TRAINING_0_DFI_RESET_N_P1_OUT ),
        .DFI_RESET_N_P2_OUT            ( IOD_TRAINING_0_DFI_RESET_N_P2_OUT ),
        .DFI_RESET_N_P3_OUT            ( IOD_TRAINING_0_DFI_RESET_N_P3_OUT ),
        .DFI_BANK_P0_OUT               ( DFI_BANK_P0_OUT_net_0 ),
        .DFI_BANK_P1_OUT               ( DFI_BANK_P1_OUT_net_0 ),
        .DFI_BANK_P2_OUT               ( DFI_BANK_P2_OUT_net_0 ),
        .DFI_BANK_P3_OUT               ( DFI_BANK_P3_OUT_net_0 ),
        .DFI_CS_N_P0_OUT               ( IOD_TRAINING_0_DFI_CS_N_P0_OUT ),
        .DFI_CS_N_P1_OUT               ( IOD_TRAINING_0_DFI_CS_N_P1_OUT ),
        .DFI_CS_N_P2_OUT               ( IOD_TRAINING_0_DFI_CS_N_P2_OUT ),
        .DFI_CS_N_P3_OUT               ( IOD_TRAINING_0_DFI_CS_N_P3_OUT ),
        .DFI_ODT_P0_OUT                ( IOD_TRAINING_0_DFI_ODT_P0_OUT ),
        .DFI_ODT_P1_OUT                ( IOD_TRAINING_0_DFI_ODT_P1_OUT ),
        .DFI_ODT_P2_OUT                ( IOD_TRAINING_0_DFI_ODT_P2_OUT ),
        .DFI_ODT_P3_OUT                ( IOD_TRAINING_0_DFI_ODT_P3_OUT ),
        .DFI_CKE_P0_OUT                ( IOD_TRAINING_0_DFI_CKE_P0_OUT ),
        .DFI_CKE_P1_OUT                ( IOD_TRAINING_0_DFI_CKE_P1_OUT ),
        .DFI_CKE_P2_OUT                ( IOD_TRAINING_0_DFI_CKE_P2_OUT ),
        .DFI_CKE_P3_OUT                ( IOD_TRAINING_0_DFI_CKE_P3_OUT ),
        .DFI_RAS_N_P0_OUT              ( IOD_TRAINING_0_DFI_RAS_N_P0_OUT ),
        .DFI_RAS_N_P1_OUT              ( IOD_TRAINING_0_DFI_RAS_N_P1_OUT ),
        .DFI_RAS_N_P2_OUT              ( IOD_TRAINING_0_DFI_RAS_N_P2_OUT ),
        .DFI_RAS_N_P3_OUT              ( IOD_TRAINING_0_DFI_RAS_N_P3_OUT ),
        .DFI_CAS_N_P0_OUT              ( IOD_TRAINING_0_DFI_CAS_N_P0_OUT ),
        .DFI_CAS_N_P1_OUT              ( IOD_TRAINING_0_DFI_CAS_N_P1_OUT ),
        .DFI_CAS_N_P2_OUT              ( IOD_TRAINING_0_DFI_CAS_N_P2_OUT ),
        .DFI_CAS_N_P3_OUT              ( IOD_TRAINING_0_DFI_CAS_N_P3_OUT ),
        .DFI_WE_N_P0_OUT               ( IOD_TRAINING_0_DFI_WE_N_P0_OUT ),
        .DFI_WE_N_P1_OUT               ( IOD_TRAINING_0_DFI_WE_N_P1_OUT ),
        .DFI_WE_N_P2_OUT               ( IOD_TRAINING_0_DFI_WE_N_P2_OUT ),
        .DFI_WE_N_P3_OUT               ( IOD_TRAINING_0_DFI_WE_N_P3_OUT ),
        .DFI_ACT_N_P0_OUT              ( IOD_TRAINING_0_DFI_ACT_N_P0_OUT ),
        .DFI_ACT_N_P1_OUT              ( IOD_TRAINING_0_DFI_ACT_N_P1_OUT ),
        .DFI_ACT_N_P2_OUT              ( IOD_TRAINING_0_DFI_ACT_N_P2_OUT ),
        .DFI_ACT_N_P3_OUT              ( IOD_TRAINING_0_DFI_ACT_N_P3_OUT ),
        .DFI_BG_P0_OUT                 ( DFI_BG_P0_OUT_net_0 ),
        .DFI_BG_P1_OUT                 ( DFI_BG_P1_OUT_net_0 ),
        .DFI_BG_P2_OUT                 ( DFI_BG_P2_OUT_net_0 ),
        .DFI_BG_P3_OUT                 ( DFI_BG_P3_OUT_net_0 ) 
        );

//--------PF_DDR4_SS_DDRPHY_BLK_IOD_WE_N_PF_IOD   -   Actel:SgCore:PF_IOD:1.0.218
PF_DDR4_SS_DDRPHY_BLK_IOD_WE_N_PF_IOD IOD_WE_N(
        // Inputs
        .ARST_N                    ( LANECTRL_ADDR_CMD_0_ARST_N ),
        .RX_SYNC_RST               ( LANECTRL_ADDR_CMD_0_RX_SYNC_RST ),
        .TX_SYNC_RST               ( LANECTRL_ADDR_CMD_0_TX_SYNC_RST ),
        .HS_IO_CLK                 ( HS_IO_CLK ),
        .TX_DQS_270                ( LANECTRL_ADDR_CMD_0_TX_DQS_270 ),
        .TX_DATA_0                 ( TX_DATA_0_net_12 ),
        .OE_DATA_0                 ( OE_DATA_0_const_net_11 ),
        .DELAY_LINE_MOVE_0         ( IOD_TRAINING_0_CMD_DELAY_LINE_MOVE ),
        .DELAY_LINE_DIRECTION_0    ( IOD_TRAINING_0_CMD_DELAY_LINE_DIRECTION ),
        .DELAY_LINE_LOAD_0         ( IOD_TRAINING_0_CMD_DELAY_LINE_LOAD ),
        .FAB_CLK                   ( SYS_CLK ),
        .ODT_EN_0                  ( GND_net ), // tied to 1'b0 from definition
        // Outputs
        .DELAY_LINE_OUT_OF_RANGE_0 (  ),
        .PAD_O                     ( WE_N_net_0 ) 
        );

//--------PF_DDR4_SS_DDRPHY_BLK_LANE_0_CTRL_PF_LANECTRL   -   Actel:SgCore:PF_LANECTRL:2.0.102
PF_DDR4_SS_DDRPHY_BLK_LANE_0_CTRL_PF_LANECTRL LANE_0_CTRL(
        // Inputs
        .DQS                        ( LANE_0_IOD_DQS_DQS ),
        .HS_IO_CLK                  ( HS_IO_CLK_net_0 ),
        .DLL_CODE                   ( DLL_CODE ),
        .FAB_CLK                    ( SYS_CLK ),
        .RESET                      ( SYNC_SYS_RST_N_net_0 ),
        .DDR_READ                   ( DFI_RDLVL_GATE_EN ),
        .READ_CLK_SEL               ( READ_CLK_SEL_net_0 ),
        .DELAY_LINE_SEL             ( IOD_TRAINING_0_DELAY_LINE_SEL_RD0to0 ),
        .DELAY_LINE_LOAD            ( IOD_TRAINING_0_LOAD8to8 ),
        .DELAY_LINE_DIRECTION       ( IOD_TRAINING_0_DIRECTION8to8 ),
        .DELAY_LINE_MOVE            ( IOD_TRAINING_0_MOVE8to8 ),
        .HS_IO_CLK_PAUSE            ( IOD_TRAINING_0_INIT_PAUSE0to0 ),
        .EYE_MONITOR_WIDTH_IN       ( EYE_MONITOR_WIDTH_IN_const_net_0 ),
        .ODT_EN                     ( VCC_net ),
        .CDR_CLK_A_SEL              ( IOD_TRAINING_0_DQSW_SELA7to0 ),
        .DDR_DO_READ                ( LANE_0_IOD_READ_TRAINING_DDR_DO_READ ),
        .SWITCH                     ( LANE_0_IOD_READ_TRAINING_SWITCH ),
        // Outputs
        .EYE_MONITOR_WIDTH_OUT      ( LANE_0_CTRL_EYE_MONITOR_WIDTH_OUT ),
        .ODT_EN_SEL                 (  ),
        .RX_DQS_90                  ( LANE_0_CTRL_RX_DQS_90 ),
        .TX_DQS                     ( LANE_0_CTRL_TX_DQS ),
        .TX_DQS_270                 ( LANE_0_CTRL_TX_DQS_270 ),
        .FIFO_WR_PTR                ( LANE_0_CTRL_FIFO_WR_PTR ),
        .FIFO_RD_PTR                ( LANE_0_CTRL_FIFO_RD_PTR ),
        .ARST_N                     ( LANE_0_CTRL_ARST_N ),
        .RX_SYNC_RST                ( LANE_0_CTRL_RX_SYNC_RST ),
        .TX_SYNC_RST                ( LANE_0_CTRL_TX_SYNC_RST ),
        .ODT_EN_OUT                 (  ),
        .RX_DATA_VALID              ( LANE_0_CTRL_RX_DATA_VALID ),
        .RX_BURST_DETECT            ( LANE_0_CTRL_RX_BURST_DETECT ),
        .RX_DELAY_LINE_OUT_OF_RANGE ( LANE_0_CTRL_RX_DELAY_LINE_OUT_OF_RANGE ),
        .TX_DELAY_LINE_OUT_OF_RANGE ( LANE_0_CTRL_TX_DELAY_LINE_OUT_OF_RANGE ),
        .A_OUT_RST_N                (  ) 
        );

//--------PF_DDR4_SS_DDRPHY_BLK_LANE_0_IOD_DM_PF_IOD   -   Actel:SgCore:PF_IOD:1.0.218
PF_DDR4_SS_DDRPHY_BLK_LANE_0_IOD_DM_PF_IOD LANE_0_IOD_DM(
        // Inputs
        .ARST_N                    ( LANE_0_CTRL_ARST_N ),
        .RX_SYNC_RST               ( LANE_0_CTRL_RX_SYNC_RST ),
        .TX_SYNC_RST               ( LANE_0_CTRL_TX_SYNC_RST ),
        .HS_IO_CLK                 ( HS_IO_CLK ),
        .TX_DQS                    ( LANE_0_CTRL_TX_DQS ),
        .TX_DATA_0                 ( TX_DATA_0_net_13 ),
        .OE_DATA_0                 ( OE_DATA_0_net_1 ),
        .DELAY_LINE_MOVE_0         ( GND_net ),
        .DELAY_LINE_DIRECTION_0    ( GND_net ),
        .DELAY_LINE_LOAD_0         ( GND_net ),
        .FAB_CLK                   ( SYS_CLK ),
        .ODT_EN_0                  ( GND_net ), // tied to 1'b0 from definition
        // Outputs
        .DELAY_LINE_OUT_OF_RANGE_0 (  ),
        .PAD_O                     ( DM_N_net_0 ),
        .RX_FB                     ( LANE_0_IOD_DM_RX_FB ) 
        );

//--------PF_DDR4_SS_DDRPHY_BLK_LANE_0_IOD_DQ_PF_IOD   -   Actel:SgCore:PF_IOD:1.0.218
PF_DDR4_SS_DDRPHY_BLK_LANE_0_IOD_DQ_PF_IOD LANE_0_IOD_DQ(
        // Inputs
        .ARST_N                    ( LANE_0_CTRL_ARST_N ),
        .RX_SYNC_RST               ( LANE_0_CTRL_RX_SYNC_RST ),
        .TX_SYNC_RST               ( LANE_0_CTRL_TX_SYNC_RST ),
        .HS_IO_CLK                 ( HS_IO_CLK ),
        .RX_DQS_90                 ( LANE_0_CTRL_RX_DQS_90 ),
        .TX_DQS                    ( LANE_0_CTRL_TX_DQS ),
        .FIFO_WR_PTR               ( LANE_0_CTRL_FIFO_WR_PTR ),
        .FIFO_RD_PTR               ( LANE_0_CTRL_FIFO_RD_PTR ),
        .EYE_MONITOR_LANE_WIDTH    ( LANE_0_CTRL_EYE_MONITOR_WIDTH_OUT ),
        .TX_DATA_0                 ( TX_DATA_0_net_14 ),
        .TX_DATA_1                 ( TX_DATA_1_net_3 ),
        .TX_DATA_2                 ( TX_DATA_2_net_1 ),
        .TX_DATA_3                 ( TX_DATA_3_net_1 ),
        .TX_DATA_4                 ( TX_DATA_4_net_1 ),
        .TX_DATA_5                 ( TX_DATA_5_net_1 ),
        .TX_DATA_6                 ( TX_DATA_6_net_1 ),
        .TX_DATA_7                 ( TX_DATA_7_net_1 ),
        .OE_DATA_0                 ( OE_DATA_0_net_2 ),
        .OE_DATA_1                 ( OE_DATA_1_net_0 ),
        .OE_DATA_2                 ( OE_DATA_2_net_0 ),
        .OE_DATA_3                 ( OE_DATA_3_net_0 ),
        .OE_DATA_4                 ( OE_DATA_4_net_0 ),
        .OE_DATA_5                 ( OE_DATA_5_net_0 ),
        .OE_DATA_6                 ( OE_DATA_6_net_0 ),
        .OE_DATA_7                 ( OE_DATA_7_net_0 ),
        .EYE_MONITOR_CLEAR_FLAGS_0 ( GND_net ),
        .EYE_MONITOR_CLEAR_FLAGS_1 ( GND_net ),
        .EYE_MONITOR_CLEAR_FLAGS_2 ( GND_net ),
        .EYE_MONITOR_CLEAR_FLAGS_3 ( GND_net ),
        .EYE_MONITOR_CLEAR_FLAGS_4 ( GND_net ),
        .EYE_MONITOR_CLEAR_FLAGS_5 ( GND_net ),
        .EYE_MONITOR_CLEAR_FLAGS_6 ( GND_net ),
        .EYE_MONITOR_CLEAR_FLAGS_7 ( GND_net ),
        .DELAY_LINE_MOVE_0         ( IOD_TRAINING_0_MOVE0to0 ),
        .DELAY_LINE_MOVE_1         ( IOD_TRAINING_0_MOVE1to1 ),
        .DELAY_LINE_MOVE_2         ( IOD_TRAINING_0_MOVE2to2 ),
        .DELAY_LINE_MOVE_3         ( IOD_TRAINING_0_MOVE3to3 ),
        .DELAY_LINE_MOVE_4         ( IOD_TRAINING_0_MOVE4to4 ),
        .DELAY_LINE_MOVE_5         ( IOD_TRAINING_0_MOVE5to5 ),
        .DELAY_LINE_MOVE_6         ( IOD_TRAINING_0_MOVE6to6 ),
        .DELAY_LINE_MOVE_7         ( IOD_TRAINING_0_MOVE7to7 ),
        .DELAY_LINE_DIRECTION_0    ( IOD_TRAINING_0_DIRECTION0to0 ),
        .DELAY_LINE_DIRECTION_1    ( IOD_TRAINING_0_DIRECTION1to1 ),
        .DELAY_LINE_DIRECTION_2    ( IOD_TRAINING_0_DIRECTION2to2 ),
        .DELAY_LINE_DIRECTION_3    ( IOD_TRAINING_0_DIRECTION3to3 ),
        .DELAY_LINE_DIRECTION_4    ( IOD_TRAINING_0_DIRECTION4to4 ),
        .DELAY_LINE_DIRECTION_5    ( IOD_TRAINING_0_DIRECTION5to5 ),
        .DELAY_LINE_DIRECTION_6    ( IOD_TRAINING_0_DIRECTION6to6 ),
        .DELAY_LINE_DIRECTION_7    ( IOD_TRAINING_0_DIRECTION7to7 ),
        .DELAY_LINE_LOAD_0         ( IOD_TRAINING_0_LOAD0to0 ),
        .DELAY_LINE_LOAD_1         ( IOD_TRAINING_0_LOAD1to1 ),
        .DELAY_LINE_LOAD_2         ( IOD_TRAINING_0_LOAD2to2 ),
        .DELAY_LINE_LOAD_3         ( IOD_TRAINING_0_LOAD3to3 ),
        .DELAY_LINE_LOAD_4         ( IOD_TRAINING_0_LOAD4to4 ),
        .DELAY_LINE_LOAD_5         ( IOD_TRAINING_0_LOAD5to5 ),
        .DELAY_LINE_LOAD_6         ( IOD_TRAINING_0_LOAD6to6 ),
        .DELAY_LINE_LOAD_7         ( IOD_TRAINING_0_LOAD7to7 ),
        .FAB_CLK                   ( SYS_CLK ),
        .ODT_EN_0                  ( GND_net ), // tied to 1'b0 from definition
        .ODT_EN_1                  ( GND_net ), // tied to 1'b0 from definition
        .ODT_EN_2                  ( GND_net ), // tied to 1'b0 from definition
        .ODT_EN_3                  ( GND_net ), // tied to 1'b0 from definition
        .ODT_EN_4                  ( GND_net ), // tied to 1'b0 from definition
        .ODT_EN_5                  ( GND_net ), // tied to 1'b0 from definition
        .ODT_EN_6                  ( GND_net ), // tied to 1'b0 from definition
        .ODT_EN_7                  ( GND_net ), // tied to 1'b0 from definition
        // Outputs
        .DELAY_LINE_OUT_OF_RANGE_0 ( LANE_0_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_0 ),
        .DELAY_LINE_OUT_OF_RANGE_1 ( LANE_0_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_1 ),
        .DELAY_LINE_OUT_OF_RANGE_2 ( LANE_0_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_2 ),
        .DELAY_LINE_OUT_OF_RANGE_3 ( LANE_0_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_3 ),
        .DELAY_LINE_OUT_OF_RANGE_4 ( LANE_0_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_4 ),
        .DELAY_LINE_OUT_OF_RANGE_5 ( LANE_0_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_5 ),
        .DELAY_LINE_OUT_OF_RANGE_6 ( LANE_0_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_6 ),
        .DELAY_LINE_OUT_OF_RANGE_7 ( LANE_0_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_7 ),
        .EYE_MONITOR_EARLY_0       (  ),
        .EYE_MONITOR_EARLY_1       (  ),
        .EYE_MONITOR_EARLY_2       (  ),
        .EYE_MONITOR_EARLY_3       (  ),
        .EYE_MONITOR_EARLY_4       (  ),
        .EYE_MONITOR_EARLY_5       (  ),
        .EYE_MONITOR_EARLY_6       (  ),
        .EYE_MONITOR_EARLY_7       (  ),
        .EYE_MONITOR_LATE_0        (  ),
        .EYE_MONITOR_LATE_1        (  ),
        .EYE_MONITOR_LATE_2        (  ),
        .EYE_MONITOR_LATE_3        (  ),
        .EYE_MONITOR_LATE_4        (  ),
        .EYE_MONITOR_LATE_5        (  ),
        .EYE_MONITOR_LATE_6        (  ),
        .EYE_MONITOR_LATE_7        (  ),
        .RX_DATA_0                 ( RX_DATA_0_net_3 ),
        .RX_DATA_1                 ( RX_DATA_1_net_0 ),
        .RX_DATA_2                 ( RX_DATA_2_net_0 ),
        .RX_DATA_3                 ( RX_DATA_3_net_0 ),
        .RX_DATA_4                 ( RX_DATA_4_net_0 ),
        .RX_DATA_5                 ( RX_DATA_5_net_0 ),
        .RX_DATA_6                 ( RX_DATA_6_net_0 ),
        .RX_DATA_7                 ( RX_DATA_7_net_0 ),
        .RX_BYPASS_DATA_0          ( LANE_0_IOD_DQ_RX_BYPASS_DATA_0 ),
        .RX_BYPASS_DATA_1          ( LANE_0_IOD_DQ_RX_BYPASS_DATA_1 ),
        .RX_BYPASS_DATA_2          ( LANE_0_IOD_DQ_RX_BYPASS_DATA_2 ),
        .RX_BYPASS_DATA_3          ( LANE_0_IOD_DQ_RX_BYPASS_DATA_3 ),
        .RX_BYPASS_DATA_4          ( LANE_0_IOD_DQ_RX_BYPASS_DATA_4 ),
        .RX_BYPASS_DATA_5          ( LANE_0_IOD_DQ_RX_BYPASS_DATA_5 ),
        .RX_BYPASS_DATA_6          ( LANE_0_IOD_DQ_RX_BYPASS_DATA_6 ),
        .RX_BYPASS_DATA_7          ( LANE_0_IOD_DQ_RX_BYPASS_DATA_7 ),
        // Inouts
        .PAD                       ( { DQ[7:7] , DQ[6:6] , DQ[5:5] , DQ[4:4] , DQ[3:3] , DQ[2:2] , DQ[1:1] , DQ[0:0] } ) 
        );

//--------PF_DDR4_SS_DDRPHY_BLK_LANE_0_IOD_DQS_PF_IOD   -   Actel:SgCore:PF_IOD:1.0.218
PF_DDR4_SS_DDRPHY_BLK_LANE_0_IOD_DQS_PF_IOD LANE_0_IOD_DQS(
        // Inputs
        .ARST_N                    ( LANE_0_CTRL_ARST_N ),
        .RX_SYNC_RST               ( LANE_0_CTRL_RX_SYNC_RST ),
        .TX_SYNC_RST               ( LANE_0_CTRL_TX_SYNC_RST ),
        .HS_IO_CLK                 ( HS_IO_CLK ),
        .RX_DQS_90                 ( LANE_0_CTRL_RX_DQS_90 ),
        .TX_DQS_270                ( LANE_0_CTRL_TX_DQS_270 ),
        .FIFO_WR_PTR               ( LANE_0_CTRL_FIFO_WR_PTR ),
        .FIFO_RD_PTR               ( LANE_0_CTRL_FIFO_RD_PTR ),
        .EYE_MONITOR_LANE_WIDTH    ( LANE_0_CTRL_EYE_MONITOR_WIDTH_OUT ),
        .TX_DATA_0                 ( TX_DATA_0_const_net_0 ),
        .OE_DATA_0                 ( OE_DATA_0_net_3 ),
        .EYE_MONITOR_CLEAR_FLAGS_0 ( GND_net ),
        .DELAY_LINE_MOVE_0         ( GND_net ),
        .DELAY_LINE_DIRECTION_0    ( GND_net ),
        .DELAY_LINE_LOAD_0         ( GND_net ),
        .FAB_CLK                   ( SYS_CLK ),
        .ODT_EN_0                  ( GND_net ), // tied to 1'b0 from definition
        // Outputs
        .DELAY_LINE_OUT_OF_RANGE_0 (  ),
        .EYE_MONITOR_EARLY_0       (  ),
        .EYE_MONITOR_LATE_0        (  ),
        .RX_DATA_0                 (  ),
        .DQS                       ( LANE_0_IOD_DQS_DQS ),
        .DQS_N                     ( LANE_0_IOD_DQS_DQS_N ),
        // Inouts
        .PAD                       ( DQS[0:0] ),
        .PAD_N                     ( DQS_N[0:0] ) 
        );

//--------PF_DDR4_SS_DDRPHY_BLK_LANE_0_IOD_DQSW_TRAINING_PF_IOD   -   Actel:SgCore:PF_IOD:1.0.218
PF_DDR4_SS_DDRPHY_BLK_LANE_0_IOD_DQSW_TRAINING_PF_IOD LANE_0_IOD_DQSW_TRAINING(
        // Inputs
        .RX_N_0                    ( LANE_0_IOD_DM_RX_FB ),
        .HS_IO_CLK                 ( HS_IO_CLK ),
        .TX_DATA_0                 ( TX_DATA_0_const_net_1 ),
        .OE_DATA_0                 ( OE_DATA_0_const_net_12 ),
        .EYE_MONITOR_CLEAR_FLAGS_0 ( IOD_TRAINING_0_DQSW_EYE_MONITOR_CLR_FLAGS0to0 ),
        .DELAY_LINE_MOVE_0         ( IOD_TRAINING_0_DQSW_DELAY_LINE_MOVE0to0 ),
        .DELAY_LINE_DIRECTION_0    ( IOD_TRAINING_0_DQSW_DELAY_LINE_DIRECTION0to0 ),
        .DELAY_LINE_LOAD_0         ( IOD_TRAINING_0_DQSW_DELAY_LINE_LOAD0to0 ),
        .FAB_CLK                   ( SYS_CLK ),
        .ODT_EN_0                  ( GND_net ), // tied to 1'b0 from definition
        // Outputs
        .TX_0                      ( LANE_0_IOD_DQSW_TRAINING_TX_0 ),
        .OE_0                      ( LANE_0_IOD_DQSW_TRAINING_OE_0 ),
        .DELAY_LINE_OUT_OF_RANGE_0 ( LANE_0_IOD_DQSW_TRAINING_DELAY_LINE_OUT_OF_RANGE_0 ),
        .EYE_MONITOR_EARLY_0       ( LANE_0_IOD_DQSW_TRAINING_EYE_MONITOR_EARLY_0 ),
        .EYE_MONITOR_LATE_0        ( LANE_0_IOD_DQSW_TRAINING_EYE_MONITOR_LATE_0 ),
        .RX_DATA_0                 ( RX_DATA_0_net_4 ) 
        );

//--------PF_DDR4_SS_DDRPHY_BLK_LANE_0_IOD_READ_TRAINING_PF_IOD   -   Actel:SgCore:PF_IOD:1.0.218
PF_DDR4_SS_DDRPHY_BLK_LANE_0_IOD_READ_TRAINING_PF_IOD LANE_0_IOD_READ_TRAINING(
        // Inputs
        .RX_P_0                    ( LANE_0_IOD_DQS_DQS_N ),
        .ARST_N                    ( LANE_0_CTRL_ARST_N ),
        .RX_SYNC_RST               ( LANE_0_CTRL_RX_SYNC_RST ),
        .TX_SYNC_RST               ( LANE_0_CTRL_TX_SYNC_RST ),
        .HS_IO_CLK                 ( HS_IO_CLK ),
        .TX_DQS                    ( LANE_0_CTRL_TX_DQS ),
        .FIFO_WR_PTR               ( LANE_0_CTRL_FIFO_WR_PTR ),
        .FIFO_RD_PTR               ( LANE_0_CTRL_FIFO_RD_PTR ),
        .TX_DATA_0                 ( TX_DATA_0_net_15 ),
        .OE_DATA_0                 ( OE_DATA_0_net_4 ),
        .EYE_MONITOR_CLEAR_FLAGS_0 ( IOD_TRAINING_0_DQSW270_EYE_MONITOR_CLR_FLAGS0to0 ),
        .DELAY_LINE_MOVE_0         ( IOD_TRAINING_0_DQSW270_DELAY_LINE_MOVE0to0 ),
        .DELAY_LINE_DIRECTION_0    ( IOD_TRAINING_0_DQSW270_DELAY_LINE_DIRECTION0to0 ),
        .DELAY_LINE_LOAD_0         ( IOD_TRAINING_0_DQSW270_DELAY_LINE_LOAD0to0 ),
        .FAB_CLK                   ( SYS_CLK ),
        .ODT_EN_0                  ( GND_net ), // tied to 1'b0 from definition
        // Outputs
        .DELAY_LINE_OUT_OF_RANGE_0 ( LANE_0_IOD_READ_TRAINING_DELAY_LINE_OUT_OF_RANGE_0 ),
        .EYE_MONITOR_EARLY_0       ( LANE_0_IOD_READ_TRAINING_EYE_MONITOR_EARLY_0 ),
        .EYE_MONITOR_LATE_0        ( LANE_0_IOD_READ_TRAINING_EYE_MONITOR_LATE_0 ),
        .RX_DATA_0                 ( RX_DATA_0_net_5 ),
        .DDR_DO_READ               ( LANE_0_IOD_READ_TRAINING_DDR_DO_READ ),
        .SWITCH                    ( LANE_0_IOD_READ_TRAINING_SWITCH ) 
        );

//--------PF_DDR4_SS_DDRPHY_BLK_LANE_1_CTRL_PF_LANECTRL   -   Actel:SgCore:PF_LANECTRL:2.0.102
PF_DDR4_SS_DDRPHY_BLK_LANE_1_CTRL_PF_LANECTRL LANE_1_CTRL(
        // Inputs
        .DQS                        ( LANE_1_IOD_DQS_DQS ),
        .HS_IO_CLK                  ( HS_IO_CLK_net_1 ),
        .DLL_CODE                   ( DLL_CODE ),
        .FAB_CLK                    ( SYS_CLK ),
        .RESET                      ( SYNC_SYS_RST_N_net_0 ),
        .DDR_READ                   ( DFI_RDLVL_GATE_EN ),
        .READ_CLK_SEL               ( READ_CLK_SEL_net_1 ),
        .DELAY_LINE_SEL             ( IOD_TRAINING_0_DELAY_LINE_SEL_RD1to1 ),
        .DELAY_LINE_LOAD            ( IOD_TRAINING_0_LOAD17to17 ),
        .DELAY_LINE_DIRECTION       ( IOD_TRAINING_0_DIRECTION17to17 ),
        .DELAY_LINE_MOVE            ( IOD_TRAINING_0_MOVE17to17 ),
        .HS_IO_CLK_PAUSE            ( IOD_TRAINING_0_INIT_PAUSE1to1 ),
        .EYE_MONITOR_WIDTH_IN       ( EYE_MONITOR_WIDTH_IN_const_net_1 ),
        .ODT_EN                     ( VCC_net ),
        .CDR_CLK_A_SEL              ( IOD_TRAINING_0_DQSW_SELA15to8 ),
        .DDR_DO_READ                ( LANE_1_IOD_READ_TRAINING_DDR_DO_READ ),
        .SWITCH                     ( LANE_1_IOD_READ_TRAINING_SWITCH ),
        // Outputs
        .EYE_MONITOR_WIDTH_OUT      ( LANE_1_CTRL_EYE_MONITOR_WIDTH_OUT ),
        .ODT_EN_SEL                 (  ),
        .RX_DQS_90                  ( LANE_1_CTRL_RX_DQS_90 ),
        .TX_DQS                     ( LANE_1_CTRL_TX_DQS ),
        .TX_DQS_270                 ( LANE_1_CTRL_TX_DQS_270 ),
        .FIFO_WR_PTR                ( LANE_1_CTRL_FIFO_WR_PTR ),
        .FIFO_RD_PTR                ( LANE_1_CTRL_FIFO_RD_PTR ),
        .ARST_N                     ( LANE_1_CTRL_ARST_N ),
        .RX_SYNC_RST                ( LANE_1_CTRL_RX_SYNC_RST ),
        .TX_SYNC_RST                ( LANE_1_CTRL_TX_SYNC_RST ),
        .ODT_EN_OUT                 (  ),
        .RX_DATA_VALID              ( LANE_1_CTRL_RX_DATA_VALID ),
        .RX_BURST_DETECT            ( LANE_1_CTRL_RX_BURST_DETECT ),
        .RX_DELAY_LINE_OUT_OF_RANGE ( LANE_1_CTRL_RX_DELAY_LINE_OUT_OF_RANGE ),
        .TX_DELAY_LINE_OUT_OF_RANGE ( LANE_1_CTRL_TX_DELAY_LINE_OUT_OF_RANGE ),
        .A_OUT_RST_N                (  ) 
        );

//--------PF_DDR4_SS_DDRPHY_BLK_LANE_1_IOD_DM_PF_IOD   -   Actel:SgCore:PF_IOD:1.0.218
PF_DDR4_SS_DDRPHY_BLK_LANE_1_IOD_DM_PF_IOD LANE_1_IOD_DM(
        // Inputs
        .ARST_N                    ( LANE_1_CTRL_ARST_N ),
        .RX_SYNC_RST               ( LANE_1_CTRL_RX_SYNC_RST ),
        .TX_SYNC_RST               ( LANE_1_CTRL_TX_SYNC_RST ),
        .HS_IO_CLK                 ( HS_IO_CLK ),
        .TX_DQS                    ( LANE_1_CTRL_TX_DQS ),
        .TX_DATA_0                 ( TX_DATA_0_net_16 ),
        .OE_DATA_0                 ( OE_DATA_0_net_5 ),
        .DELAY_LINE_MOVE_0         ( GND_net ),
        .DELAY_LINE_DIRECTION_0    ( GND_net ),
        .DELAY_LINE_LOAD_0         ( GND_net ),
        .FAB_CLK                   ( SYS_CLK ),
        .ODT_EN_0                  ( GND_net ), // tied to 1'b0 from definition
        // Outputs
        .DELAY_LINE_OUT_OF_RANGE_0 (  ),
        .PAD_O                     ( DM_N_0 ),
        .RX_FB                     ( LANE_1_IOD_DM_RX_FB ) 
        );

//--------PF_DDR4_SS_DDRPHY_BLK_LANE_1_IOD_DQ_PF_IOD   -   Actel:SgCore:PF_IOD:1.0.218
PF_DDR4_SS_DDRPHY_BLK_LANE_1_IOD_DQ_PF_IOD LANE_1_IOD_DQ(
        // Inputs
        .ARST_N                    ( LANE_1_CTRL_ARST_N ),
        .RX_SYNC_RST               ( LANE_1_CTRL_RX_SYNC_RST ),
        .TX_SYNC_RST               ( LANE_1_CTRL_TX_SYNC_RST ),
        .HS_IO_CLK                 ( HS_IO_CLK ),
        .RX_DQS_90                 ( LANE_1_CTRL_RX_DQS_90 ),
        .TX_DQS                    ( LANE_1_CTRL_TX_DQS ),
        .FIFO_WR_PTR               ( LANE_1_CTRL_FIFO_WR_PTR ),
        .FIFO_RD_PTR               ( LANE_1_CTRL_FIFO_RD_PTR ),
        .EYE_MONITOR_LANE_WIDTH    ( LANE_1_CTRL_EYE_MONITOR_WIDTH_OUT ),
        .TX_DATA_0                 ( TX_DATA_0_net_17 ),
        .TX_DATA_1                 ( TX_DATA_1_net_4 ),
        .TX_DATA_2                 ( TX_DATA_2_net_2 ),
        .TX_DATA_3                 ( TX_DATA_3_net_2 ),
        .TX_DATA_4                 ( TX_DATA_4_net_2 ),
        .TX_DATA_5                 ( TX_DATA_5_net_2 ),
        .TX_DATA_6                 ( TX_DATA_6_net_2 ),
        .TX_DATA_7                 ( TX_DATA_7_net_2 ),
        .OE_DATA_0                 ( OE_DATA_0_net_6 ),
        .OE_DATA_1                 ( OE_DATA_1_net_1 ),
        .OE_DATA_2                 ( OE_DATA_2_net_1 ),
        .OE_DATA_3                 ( OE_DATA_3_net_1 ),
        .OE_DATA_4                 ( OE_DATA_4_net_1 ),
        .OE_DATA_5                 ( OE_DATA_5_net_1 ),
        .OE_DATA_6                 ( OE_DATA_6_net_1 ),
        .OE_DATA_7                 ( OE_DATA_7_net_1 ),
        .EYE_MONITOR_CLEAR_FLAGS_0 ( GND_net ),
        .EYE_MONITOR_CLEAR_FLAGS_1 ( GND_net ),
        .EYE_MONITOR_CLEAR_FLAGS_2 ( GND_net ),
        .EYE_MONITOR_CLEAR_FLAGS_3 ( GND_net ),
        .EYE_MONITOR_CLEAR_FLAGS_4 ( GND_net ),
        .EYE_MONITOR_CLEAR_FLAGS_5 ( GND_net ),
        .EYE_MONITOR_CLEAR_FLAGS_6 ( GND_net ),
        .EYE_MONITOR_CLEAR_FLAGS_7 ( GND_net ),
        .DELAY_LINE_MOVE_0         ( IOD_TRAINING_0_MOVE9to9 ),
        .DELAY_LINE_MOVE_1         ( IOD_TRAINING_0_MOVE10to10 ),
        .DELAY_LINE_MOVE_2         ( IOD_TRAINING_0_MOVE11to11 ),
        .DELAY_LINE_MOVE_3         ( IOD_TRAINING_0_MOVE12to12 ),
        .DELAY_LINE_MOVE_4         ( IOD_TRAINING_0_MOVE13to13 ),
        .DELAY_LINE_MOVE_5         ( IOD_TRAINING_0_MOVE14to14 ),
        .DELAY_LINE_MOVE_6         ( IOD_TRAINING_0_MOVE15to15 ),
        .DELAY_LINE_MOVE_7         ( IOD_TRAINING_0_MOVE16to16 ),
        .DELAY_LINE_DIRECTION_0    ( IOD_TRAINING_0_DIRECTION9to9 ),
        .DELAY_LINE_DIRECTION_1    ( IOD_TRAINING_0_DIRECTION10to10 ),
        .DELAY_LINE_DIRECTION_2    ( IOD_TRAINING_0_DIRECTION11to11 ),
        .DELAY_LINE_DIRECTION_3    ( IOD_TRAINING_0_DIRECTION12to12 ),
        .DELAY_LINE_DIRECTION_4    ( IOD_TRAINING_0_DIRECTION13to13 ),
        .DELAY_LINE_DIRECTION_5    ( IOD_TRAINING_0_DIRECTION14to14 ),
        .DELAY_LINE_DIRECTION_6    ( IOD_TRAINING_0_DIRECTION15to15 ),
        .DELAY_LINE_DIRECTION_7    ( IOD_TRAINING_0_DIRECTION16to16 ),
        .DELAY_LINE_LOAD_0         ( IOD_TRAINING_0_LOAD9to9 ),
        .DELAY_LINE_LOAD_1         ( IOD_TRAINING_0_LOAD10to10 ),
        .DELAY_LINE_LOAD_2         ( IOD_TRAINING_0_LOAD11to11 ),
        .DELAY_LINE_LOAD_3         ( IOD_TRAINING_0_LOAD12to12 ),
        .DELAY_LINE_LOAD_4         ( IOD_TRAINING_0_LOAD13to13 ),
        .DELAY_LINE_LOAD_5         ( IOD_TRAINING_0_LOAD14to14 ),
        .DELAY_LINE_LOAD_6         ( IOD_TRAINING_0_LOAD15to15 ),
        .DELAY_LINE_LOAD_7         ( IOD_TRAINING_0_LOAD16to16 ),
        .FAB_CLK                   ( SYS_CLK ),
        .ODT_EN_0                  ( GND_net ), // tied to 1'b0 from definition
        .ODT_EN_1                  ( GND_net ), // tied to 1'b0 from definition
        .ODT_EN_2                  ( GND_net ), // tied to 1'b0 from definition
        .ODT_EN_3                  ( GND_net ), // tied to 1'b0 from definition
        .ODT_EN_4                  ( GND_net ), // tied to 1'b0 from definition
        .ODT_EN_5                  ( GND_net ), // tied to 1'b0 from definition
        .ODT_EN_6                  ( GND_net ), // tied to 1'b0 from definition
        .ODT_EN_7                  ( GND_net ), // tied to 1'b0 from definition
        // Outputs
        .DELAY_LINE_OUT_OF_RANGE_0 ( LANE_1_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_0 ),
        .DELAY_LINE_OUT_OF_RANGE_1 ( LANE_1_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_1 ),
        .DELAY_LINE_OUT_OF_RANGE_2 ( LANE_1_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_2 ),
        .DELAY_LINE_OUT_OF_RANGE_3 ( LANE_1_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_3 ),
        .DELAY_LINE_OUT_OF_RANGE_4 ( LANE_1_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_4 ),
        .DELAY_LINE_OUT_OF_RANGE_5 ( LANE_1_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_5 ),
        .DELAY_LINE_OUT_OF_RANGE_6 ( LANE_1_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_6 ),
        .DELAY_LINE_OUT_OF_RANGE_7 ( LANE_1_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_7 ),
        .EYE_MONITOR_EARLY_0       (  ),
        .EYE_MONITOR_EARLY_1       (  ),
        .EYE_MONITOR_EARLY_2       (  ),
        .EYE_MONITOR_EARLY_3       (  ),
        .EYE_MONITOR_EARLY_4       (  ),
        .EYE_MONITOR_EARLY_5       (  ),
        .EYE_MONITOR_EARLY_6       (  ),
        .EYE_MONITOR_EARLY_7       (  ),
        .EYE_MONITOR_LATE_0        (  ),
        .EYE_MONITOR_LATE_1        (  ),
        .EYE_MONITOR_LATE_2        (  ),
        .EYE_MONITOR_LATE_3        (  ),
        .EYE_MONITOR_LATE_4        (  ),
        .EYE_MONITOR_LATE_5        (  ),
        .EYE_MONITOR_LATE_6        (  ),
        .EYE_MONITOR_LATE_7        (  ),
        .RX_DATA_0                 ( RX_DATA_0_net_6 ),
        .RX_DATA_1                 ( RX_DATA_1_net_1 ),
        .RX_DATA_2                 ( RX_DATA_2_net_1 ),
        .RX_DATA_3                 ( RX_DATA_3_net_1 ),
        .RX_DATA_4                 ( RX_DATA_4_net_1 ),
        .RX_DATA_5                 ( RX_DATA_5_net_1 ),
        .RX_DATA_6                 ( RX_DATA_6_net_1 ),
        .RX_DATA_7                 ( RX_DATA_7_net_1 ),
        .RX_BYPASS_DATA_0          ( LANE_1_IOD_DQ_RX_BYPASS_DATA_0 ),
        .RX_BYPASS_DATA_1          ( LANE_1_IOD_DQ_RX_BYPASS_DATA_1 ),
        .RX_BYPASS_DATA_2          ( LANE_1_IOD_DQ_RX_BYPASS_DATA_2 ),
        .RX_BYPASS_DATA_3          ( LANE_1_IOD_DQ_RX_BYPASS_DATA_3 ),
        .RX_BYPASS_DATA_4          ( LANE_1_IOD_DQ_RX_BYPASS_DATA_4 ),
        .RX_BYPASS_DATA_5          ( LANE_1_IOD_DQ_RX_BYPASS_DATA_5 ),
        .RX_BYPASS_DATA_6          ( LANE_1_IOD_DQ_RX_BYPASS_DATA_6 ),
        .RX_BYPASS_DATA_7          ( LANE_1_IOD_DQ_RX_BYPASS_DATA_7 ),
        // Inouts
        .PAD                       ( { DQ[15:15] , DQ[14:14] , DQ[13:13] , DQ[12:12] , DQ[11:11] , DQ[10:10] , DQ[9:9] , DQ[8:8] } ) 
        );

//--------PF_DDR4_SS_DDRPHY_BLK_LANE_1_IOD_DQS_PF_IOD   -   Actel:SgCore:PF_IOD:1.0.218
PF_DDR4_SS_DDRPHY_BLK_LANE_1_IOD_DQS_PF_IOD LANE_1_IOD_DQS(
        // Inputs
        .ARST_N                    ( LANE_1_CTRL_ARST_N ),
        .RX_SYNC_RST               ( LANE_1_CTRL_RX_SYNC_RST ),
        .TX_SYNC_RST               ( LANE_1_CTRL_TX_SYNC_RST ),
        .HS_IO_CLK                 ( HS_IO_CLK ),
        .RX_DQS_90                 ( LANE_1_CTRL_RX_DQS_90 ),
        .TX_DQS_270                ( LANE_1_CTRL_TX_DQS_270 ),
        .FIFO_WR_PTR               ( LANE_1_CTRL_FIFO_WR_PTR ),
        .FIFO_RD_PTR               ( LANE_1_CTRL_FIFO_RD_PTR ),
        .EYE_MONITOR_LANE_WIDTH    ( LANE_1_CTRL_EYE_MONITOR_WIDTH_OUT ),
        .TX_DATA_0                 ( TX_DATA_0_const_net_2 ),
        .OE_DATA_0                 ( OE_DATA_0_net_7 ),
        .EYE_MONITOR_CLEAR_FLAGS_0 ( GND_net ),
        .DELAY_LINE_MOVE_0         ( GND_net ),
        .DELAY_LINE_DIRECTION_0    ( GND_net ),
        .DELAY_LINE_LOAD_0         ( GND_net ),
        .FAB_CLK                   ( SYS_CLK ),
        .ODT_EN_0                  ( GND_net ), // tied to 1'b0 from definition
        // Outputs
        .DELAY_LINE_OUT_OF_RANGE_0 (  ),
        .EYE_MONITOR_EARLY_0       (  ),
        .EYE_MONITOR_LATE_0        (  ),
        .RX_DATA_0                 (  ),
        .DQS                       ( LANE_1_IOD_DQS_DQS ),
        .DQS_N                     ( LANE_1_IOD_DQS_DQS_N ),
        // Inouts
        .PAD                       ( DQS[1:1] ),
        .PAD_N                     ( DQS_N[1:1] ) 
        );

//--------PF_DDR4_SS_DDRPHY_BLK_LANE_1_IOD_DQSW_TRAINING_PF_IOD   -   Actel:SgCore:PF_IOD:1.0.218
PF_DDR4_SS_DDRPHY_BLK_LANE_1_IOD_DQSW_TRAINING_PF_IOD LANE_1_IOD_DQSW_TRAINING(
        // Inputs
        .RX_N_0                    ( LANE_1_IOD_DM_RX_FB ),
        .HS_IO_CLK                 ( HS_IO_CLK ),
        .TX_DATA_0                 ( TX_DATA_0_const_net_3 ),
        .OE_DATA_0                 ( OE_DATA_0_const_net_13 ),
        .EYE_MONITOR_CLEAR_FLAGS_0 ( IOD_TRAINING_0_DQSW_EYE_MONITOR_CLR_FLAGS1to1 ),
        .DELAY_LINE_MOVE_0         ( IOD_TRAINING_0_DQSW_DELAY_LINE_MOVE1to1 ),
        .DELAY_LINE_DIRECTION_0    ( IOD_TRAINING_0_DQSW_DELAY_LINE_DIRECTION1to1 ),
        .DELAY_LINE_LOAD_0         ( IOD_TRAINING_0_DQSW_DELAY_LINE_LOAD1to1 ),
        .FAB_CLK                   ( SYS_CLK ),
        .ODT_EN_0                  ( GND_net ), // tied to 1'b0 from definition
        // Outputs
        .TX_0                      ( LANE_1_IOD_DQSW_TRAINING_TX_0 ),
        .OE_0                      ( LANE_1_IOD_DQSW_TRAINING_OE_0 ),
        .DELAY_LINE_OUT_OF_RANGE_0 ( LANE_1_IOD_DQSW_TRAINING_DELAY_LINE_OUT_OF_RANGE_0 ),
        .EYE_MONITOR_EARLY_0       ( LANE_1_IOD_DQSW_TRAINING_EYE_MONITOR_EARLY_0 ),
        .EYE_MONITOR_LATE_0        ( LANE_1_IOD_DQSW_TRAINING_EYE_MONITOR_LATE_0 ),
        .RX_DATA_0                 ( RX_DATA_0_net_7 ) 
        );

//--------PF_DDR4_SS_DDRPHY_BLK_LANE_1_IOD_READ_TRAINING_PF_IOD   -   Actel:SgCore:PF_IOD:1.0.218
PF_DDR4_SS_DDRPHY_BLK_LANE_1_IOD_READ_TRAINING_PF_IOD LANE_1_IOD_READ_TRAINING(
        // Inputs
        .RX_P_0                    ( LANE_1_IOD_DQS_DQS_N ),
        .ARST_N                    ( LANE_1_CTRL_ARST_N ),
        .RX_SYNC_RST               ( LANE_1_CTRL_RX_SYNC_RST ),
        .TX_SYNC_RST               ( LANE_1_CTRL_TX_SYNC_RST ),
        .HS_IO_CLK                 ( HS_IO_CLK ),
        .TX_DQS                    ( LANE_1_CTRL_TX_DQS ),
        .FIFO_WR_PTR               ( LANE_1_CTRL_FIFO_WR_PTR ),
        .FIFO_RD_PTR               ( LANE_1_CTRL_FIFO_RD_PTR ),
        .TX_DATA_0                 ( TX_DATA_0_net_18 ),
        .OE_DATA_0                 ( OE_DATA_0_net_8 ),
        .EYE_MONITOR_CLEAR_FLAGS_0 ( IOD_TRAINING_0_DQSW270_EYE_MONITOR_CLR_FLAGS1to1 ),
        .DELAY_LINE_MOVE_0         ( IOD_TRAINING_0_DQSW270_DELAY_LINE_MOVE1to1 ),
        .DELAY_LINE_DIRECTION_0    ( IOD_TRAINING_0_DQSW270_DELAY_LINE_DIRECTION1to1 ),
        .DELAY_LINE_LOAD_0         ( IOD_TRAINING_0_DQSW270_DELAY_LINE_LOAD1to1 ),
        .FAB_CLK                   ( SYS_CLK ),
        .ODT_EN_0                  ( GND_net ), // tied to 1'b0 from definition
        // Outputs
        .DELAY_LINE_OUT_OF_RANGE_0 ( LANE_1_IOD_READ_TRAINING_DELAY_LINE_OUT_OF_RANGE_0 ),
        .EYE_MONITOR_EARLY_0       ( LANE_1_IOD_READ_TRAINING_EYE_MONITOR_EARLY_0 ),
        .EYE_MONITOR_LATE_0        ( LANE_1_IOD_READ_TRAINING_EYE_MONITOR_LATE_0 ),
        .RX_DATA_0                 ( RX_DATA_0_net_8 ),
        .DDR_DO_READ               ( LANE_1_IOD_READ_TRAINING_DDR_DO_READ ),
        .SWITCH                    ( LANE_1_IOD_READ_TRAINING_SWITCH ) 
        );

//--------PF_DDR4_SS_DDRPHY_BLK_LANE_2_CTRL_PF_LANECTRL   -   Actel:SgCore:PF_LANECTRL:2.0.102
PF_DDR4_SS_DDRPHY_BLK_LANE_2_CTRL_PF_LANECTRL LANE_2_CTRL(
        // Inputs
        .DQS                        ( LANE_2_IOD_DQS_DQS ),
        .HS_IO_CLK                  ( HS_IO_CLK_net_2 ),
        .DLL_CODE                   ( DLL_CODE ),
        .FAB_CLK                    ( SYS_CLK ),
        .RESET                      ( SYNC_SYS_RST_N_net_0 ),
        .DDR_READ                   ( DFI_RDLVL_GATE_EN ),
        .READ_CLK_SEL               ( READ_CLK_SEL_net_2 ),
        .DELAY_LINE_SEL             ( IOD_TRAINING_0_DELAY_LINE_SEL_RD2to2 ),
        .DELAY_LINE_LOAD            ( IOD_TRAINING_0_LOAD26to26 ),
        .DELAY_LINE_DIRECTION       ( IOD_TRAINING_0_DIRECTION26to26 ),
        .DELAY_LINE_MOVE            ( IOD_TRAINING_0_MOVE26to26 ),
        .HS_IO_CLK_PAUSE            ( IOD_TRAINING_0_INIT_PAUSE2to2 ),
        .EYE_MONITOR_WIDTH_IN       ( EYE_MONITOR_WIDTH_IN_const_net_2 ),
        .ODT_EN                     ( VCC_net ),
        .CDR_CLK_A_SEL              ( IOD_TRAINING_0_DQSW_SELA23to16 ),
        .DDR_DO_READ                ( LANE_2_IOD_READ_TRAINING_DDR_DO_READ ),
        .SWITCH                     ( LANE_2_IOD_READ_TRAINING_SWITCH ),
        // Outputs
        .EYE_MONITOR_WIDTH_OUT      ( LANE_2_CTRL_EYE_MONITOR_WIDTH_OUT ),
        .ODT_EN_SEL                 (  ),
        .RX_DQS_90                  ( LANE_2_CTRL_RX_DQS_90 ),
        .TX_DQS                     ( LANE_2_CTRL_TX_DQS ),
        .TX_DQS_270                 ( LANE_2_CTRL_TX_DQS_270 ),
        .FIFO_WR_PTR                ( LANE_2_CTRL_FIFO_WR_PTR ),
        .FIFO_RD_PTR                ( LANE_2_CTRL_FIFO_RD_PTR ),
        .ARST_N                     ( LANE_2_CTRL_ARST_N ),
        .RX_SYNC_RST                ( LANE_2_CTRL_RX_SYNC_RST ),
        .TX_SYNC_RST                ( LANE_2_CTRL_TX_SYNC_RST ),
        .ODT_EN_OUT                 (  ),
        .RX_DATA_VALID              ( LANE_2_CTRL_RX_DATA_VALID ),
        .RX_BURST_DETECT            ( LANE_2_CTRL_RX_BURST_DETECT ),
        .RX_DELAY_LINE_OUT_OF_RANGE ( LANE_2_CTRL_RX_DELAY_LINE_OUT_OF_RANGE ),
        .TX_DELAY_LINE_OUT_OF_RANGE ( LANE_2_CTRL_TX_DELAY_LINE_OUT_OF_RANGE ),
        .A_OUT_RST_N                (  ) 
        );

//--------PF_DDR4_SS_DDRPHY_BLK_LANE_2_IOD_DM_PF_IOD   -   Actel:SgCore:PF_IOD:1.0.218
PF_DDR4_SS_DDRPHY_BLK_LANE_2_IOD_DM_PF_IOD LANE_2_IOD_DM(
        // Inputs
        .ARST_N                    ( LANE_2_CTRL_ARST_N ),
        .RX_SYNC_RST               ( LANE_2_CTRL_RX_SYNC_RST ),
        .TX_SYNC_RST               ( LANE_2_CTRL_TX_SYNC_RST ),
        .HS_IO_CLK                 ( HS_IO_CLK ),
        .TX_DQS                    ( LANE_2_CTRL_TX_DQS ),
        .TX_DATA_0                 ( TX_DATA_0_net_19 ),
        .OE_DATA_0                 ( OE_DATA_0_net_9 ),
        .DELAY_LINE_MOVE_0         ( GND_net ),
        .DELAY_LINE_DIRECTION_0    ( GND_net ),
        .DELAY_LINE_LOAD_0         ( GND_net ),
        .FAB_CLK                   ( SYS_CLK ),
        .ODT_EN_0                  ( GND_net ), // tied to 1'b0 from definition
        // Outputs
        .DELAY_LINE_OUT_OF_RANGE_0 (  ),
        .PAD_O                     ( DM_N_1 ),
        .RX_FB                     ( LANE_2_IOD_DM_RX_FB ) 
        );

//--------PF_DDR4_SS_DDRPHY_BLK_LANE_2_IOD_DQ_PF_IOD   -   Actel:SgCore:PF_IOD:1.0.218
PF_DDR4_SS_DDRPHY_BLK_LANE_2_IOD_DQ_PF_IOD LANE_2_IOD_DQ(
        // Inputs
        .ARST_N                    ( LANE_2_CTRL_ARST_N ),
        .RX_SYNC_RST               ( LANE_2_CTRL_RX_SYNC_RST ),
        .TX_SYNC_RST               ( LANE_2_CTRL_TX_SYNC_RST ),
        .HS_IO_CLK                 ( HS_IO_CLK ),
        .RX_DQS_90                 ( LANE_2_CTRL_RX_DQS_90 ),
        .TX_DQS                    ( LANE_2_CTRL_TX_DQS ),
        .FIFO_WR_PTR               ( LANE_2_CTRL_FIFO_WR_PTR ),
        .FIFO_RD_PTR               ( LANE_2_CTRL_FIFO_RD_PTR ),
        .EYE_MONITOR_LANE_WIDTH    ( LANE_2_CTRL_EYE_MONITOR_WIDTH_OUT ),
        .TX_DATA_0                 ( TX_DATA_0_net_20 ),
        .TX_DATA_1                 ( TX_DATA_1_net_5 ),
        .TX_DATA_2                 ( TX_DATA_2_net_3 ),
        .TX_DATA_3                 ( TX_DATA_3_net_3 ),
        .TX_DATA_4                 ( TX_DATA_4_net_3 ),
        .TX_DATA_5                 ( TX_DATA_5_net_3 ),
        .TX_DATA_6                 ( TX_DATA_6_net_3 ),
        .TX_DATA_7                 ( TX_DATA_7_net_3 ),
        .OE_DATA_0                 ( OE_DATA_0_net_10 ),
        .OE_DATA_1                 ( OE_DATA_1_net_2 ),
        .OE_DATA_2                 ( OE_DATA_2_net_2 ),
        .OE_DATA_3                 ( OE_DATA_3_net_2 ),
        .OE_DATA_4                 ( OE_DATA_4_net_2 ),
        .OE_DATA_5                 ( OE_DATA_5_net_2 ),
        .OE_DATA_6                 ( OE_DATA_6_net_2 ),
        .OE_DATA_7                 ( OE_DATA_7_net_2 ),
        .EYE_MONITOR_CLEAR_FLAGS_0 ( GND_net ),
        .EYE_MONITOR_CLEAR_FLAGS_1 ( GND_net ),
        .EYE_MONITOR_CLEAR_FLAGS_2 ( GND_net ),
        .EYE_MONITOR_CLEAR_FLAGS_3 ( GND_net ),
        .EYE_MONITOR_CLEAR_FLAGS_4 ( GND_net ),
        .EYE_MONITOR_CLEAR_FLAGS_5 ( GND_net ),
        .EYE_MONITOR_CLEAR_FLAGS_6 ( GND_net ),
        .EYE_MONITOR_CLEAR_FLAGS_7 ( GND_net ),
        .DELAY_LINE_MOVE_0         ( IOD_TRAINING_0_MOVE18to18 ),
        .DELAY_LINE_MOVE_1         ( IOD_TRAINING_0_MOVE19to19 ),
        .DELAY_LINE_MOVE_2         ( IOD_TRAINING_0_MOVE20to20 ),
        .DELAY_LINE_MOVE_3         ( IOD_TRAINING_0_MOVE21to21 ),
        .DELAY_LINE_MOVE_4         ( IOD_TRAINING_0_MOVE22to22 ),
        .DELAY_LINE_MOVE_5         ( IOD_TRAINING_0_MOVE23to23 ),
        .DELAY_LINE_MOVE_6         ( IOD_TRAINING_0_MOVE24to24 ),
        .DELAY_LINE_MOVE_7         ( IOD_TRAINING_0_MOVE25to25 ),
        .DELAY_LINE_DIRECTION_0    ( IOD_TRAINING_0_DIRECTION18to18 ),
        .DELAY_LINE_DIRECTION_1    ( IOD_TRAINING_0_DIRECTION19to19 ),
        .DELAY_LINE_DIRECTION_2    ( IOD_TRAINING_0_DIRECTION20to20 ),
        .DELAY_LINE_DIRECTION_3    ( IOD_TRAINING_0_DIRECTION21to21 ),
        .DELAY_LINE_DIRECTION_4    ( IOD_TRAINING_0_DIRECTION22to22 ),
        .DELAY_LINE_DIRECTION_5    ( IOD_TRAINING_0_DIRECTION23to23 ),
        .DELAY_LINE_DIRECTION_6    ( IOD_TRAINING_0_DIRECTION24to24 ),
        .DELAY_LINE_DIRECTION_7    ( IOD_TRAINING_0_DIRECTION25to25 ),
        .DELAY_LINE_LOAD_0         ( IOD_TRAINING_0_LOAD18to18 ),
        .DELAY_LINE_LOAD_1         ( IOD_TRAINING_0_LOAD19to19 ),
        .DELAY_LINE_LOAD_2         ( IOD_TRAINING_0_LOAD20to20 ),
        .DELAY_LINE_LOAD_3         ( IOD_TRAINING_0_LOAD21to21 ),
        .DELAY_LINE_LOAD_4         ( IOD_TRAINING_0_LOAD22to22 ),
        .DELAY_LINE_LOAD_5         ( IOD_TRAINING_0_LOAD23to23 ),
        .DELAY_LINE_LOAD_6         ( IOD_TRAINING_0_LOAD24to24 ),
        .DELAY_LINE_LOAD_7         ( IOD_TRAINING_0_LOAD25to25 ),
        .FAB_CLK                   ( SYS_CLK ),
        .ODT_EN_0                  ( GND_net ), // tied to 1'b0 from definition
        .ODT_EN_1                  ( GND_net ), // tied to 1'b0 from definition
        .ODT_EN_2                  ( GND_net ), // tied to 1'b0 from definition
        .ODT_EN_3                  ( GND_net ), // tied to 1'b0 from definition
        .ODT_EN_4                  ( GND_net ), // tied to 1'b0 from definition
        .ODT_EN_5                  ( GND_net ), // tied to 1'b0 from definition
        .ODT_EN_6                  ( GND_net ), // tied to 1'b0 from definition
        .ODT_EN_7                  ( GND_net ), // tied to 1'b0 from definition
        // Outputs
        .DELAY_LINE_OUT_OF_RANGE_0 ( LANE_2_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_0 ),
        .DELAY_LINE_OUT_OF_RANGE_1 ( LANE_2_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_1 ),
        .DELAY_LINE_OUT_OF_RANGE_2 ( LANE_2_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_2 ),
        .DELAY_LINE_OUT_OF_RANGE_3 ( LANE_2_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_3 ),
        .DELAY_LINE_OUT_OF_RANGE_4 ( LANE_2_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_4 ),
        .DELAY_LINE_OUT_OF_RANGE_5 ( LANE_2_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_5 ),
        .DELAY_LINE_OUT_OF_RANGE_6 ( LANE_2_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_6 ),
        .DELAY_LINE_OUT_OF_RANGE_7 ( LANE_2_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_7 ),
        .EYE_MONITOR_EARLY_0       (  ),
        .EYE_MONITOR_EARLY_1       (  ),
        .EYE_MONITOR_EARLY_2       (  ),
        .EYE_MONITOR_EARLY_3       (  ),
        .EYE_MONITOR_EARLY_4       (  ),
        .EYE_MONITOR_EARLY_5       (  ),
        .EYE_MONITOR_EARLY_6       (  ),
        .EYE_MONITOR_EARLY_7       (  ),
        .EYE_MONITOR_LATE_0        (  ),
        .EYE_MONITOR_LATE_1        (  ),
        .EYE_MONITOR_LATE_2        (  ),
        .EYE_MONITOR_LATE_3        (  ),
        .EYE_MONITOR_LATE_4        (  ),
        .EYE_MONITOR_LATE_5        (  ),
        .EYE_MONITOR_LATE_6        (  ),
        .EYE_MONITOR_LATE_7        (  ),
        .RX_DATA_0                 ( RX_DATA_0_net_9 ),
        .RX_DATA_1                 ( RX_DATA_1_net_2 ),
        .RX_DATA_2                 ( RX_DATA_2_net_2 ),
        .RX_DATA_3                 ( RX_DATA_3_net_2 ),
        .RX_DATA_4                 ( RX_DATA_4_net_2 ),
        .RX_DATA_5                 ( RX_DATA_5_net_2 ),
        .RX_DATA_6                 ( RX_DATA_6_net_2 ),
        .RX_DATA_7                 ( RX_DATA_7_net_2 ),
        .RX_BYPASS_DATA_0          ( LANE_2_IOD_DQ_RX_BYPASS_DATA_0 ),
        .RX_BYPASS_DATA_1          ( LANE_2_IOD_DQ_RX_BYPASS_DATA_1 ),
        .RX_BYPASS_DATA_2          ( LANE_2_IOD_DQ_RX_BYPASS_DATA_2 ),
        .RX_BYPASS_DATA_3          ( LANE_2_IOD_DQ_RX_BYPASS_DATA_3 ),
        .RX_BYPASS_DATA_4          ( LANE_2_IOD_DQ_RX_BYPASS_DATA_4 ),
        .RX_BYPASS_DATA_5          ( LANE_2_IOD_DQ_RX_BYPASS_DATA_5 ),
        .RX_BYPASS_DATA_6          ( LANE_2_IOD_DQ_RX_BYPASS_DATA_6 ),
        .RX_BYPASS_DATA_7          ( LANE_2_IOD_DQ_RX_BYPASS_DATA_7 ),
        // Inouts
        .PAD                       ( { DQ[23:23] , DQ[22:22] , DQ[21:21] , DQ[20:20] , DQ[19:19] , DQ[18:18] , DQ[17:17] , DQ[16:16] } ) 
        );

//--------PF_DDR4_SS_DDRPHY_BLK_LANE_2_IOD_DQS_PF_IOD   -   Actel:SgCore:PF_IOD:1.0.218
PF_DDR4_SS_DDRPHY_BLK_LANE_2_IOD_DQS_PF_IOD LANE_2_IOD_DQS(
        // Inputs
        .ARST_N                    ( LANE_2_CTRL_ARST_N ),
        .RX_SYNC_RST               ( LANE_2_CTRL_RX_SYNC_RST ),
        .TX_SYNC_RST               ( LANE_2_CTRL_TX_SYNC_RST ),
        .HS_IO_CLK                 ( HS_IO_CLK ),
        .RX_DQS_90                 ( LANE_2_CTRL_RX_DQS_90 ),
        .TX_DQS_270                ( LANE_2_CTRL_TX_DQS_270 ),
        .FIFO_WR_PTR               ( LANE_2_CTRL_FIFO_WR_PTR ),
        .FIFO_RD_PTR               ( LANE_2_CTRL_FIFO_RD_PTR ),
        .EYE_MONITOR_LANE_WIDTH    ( LANE_2_CTRL_EYE_MONITOR_WIDTH_OUT ),
        .TX_DATA_0                 ( TX_DATA_0_const_net_4 ),
        .OE_DATA_0                 ( OE_DATA_0_net_11 ),
        .EYE_MONITOR_CLEAR_FLAGS_0 ( GND_net ),
        .DELAY_LINE_MOVE_0         ( GND_net ),
        .DELAY_LINE_DIRECTION_0    ( GND_net ),
        .DELAY_LINE_LOAD_0         ( GND_net ),
        .FAB_CLK                   ( SYS_CLK ),
        .ODT_EN_0                  ( GND_net ), // tied to 1'b0 from definition
        // Outputs
        .DELAY_LINE_OUT_OF_RANGE_0 (  ),
        .EYE_MONITOR_EARLY_0       (  ),
        .EYE_MONITOR_LATE_0        (  ),
        .RX_DATA_0                 (  ),
        .DQS                       ( LANE_2_IOD_DQS_DQS ),
        .DQS_N                     ( LANE_2_IOD_DQS_DQS_N ),
        // Inouts
        .PAD                       ( DQS[2:2] ),
        .PAD_N                     ( DQS_N[2:2] ) 
        );

//--------PF_DDR4_SS_DDRPHY_BLK_LANE_2_IOD_DQSW_TRAINING_PF_IOD   -   Actel:SgCore:PF_IOD:1.0.218
PF_DDR4_SS_DDRPHY_BLK_LANE_2_IOD_DQSW_TRAINING_PF_IOD LANE_2_IOD_DQSW_TRAINING(
        // Inputs
        .RX_N_0                    ( LANE_2_IOD_DM_RX_FB ),
        .HS_IO_CLK                 ( HS_IO_CLK ),
        .TX_DATA_0                 ( TX_DATA_0_const_net_5 ),
        .OE_DATA_0                 ( OE_DATA_0_const_net_14 ),
        .EYE_MONITOR_CLEAR_FLAGS_0 ( IOD_TRAINING_0_DQSW_EYE_MONITOR_CLR_FLAGS2to2 ),
        .DELAY_LINE_MOVE_0         ( IOD_TRAINING_0_DQSW_DELAY_LINE_MOVE2to2 ),
        .DELAY_LINE_DIRECTION_0    ( IOD_TRAINING_0_DQSW_DELAY_LINE_DIRECTION2to2 ),
        .DELAY_LINE_LOAD_0         ( IOD_TRAINING_0_DQSW_DELAY_LINE_LOAD2to2 ),
        .FAB_CLK                   ( SYS_CLK ),
        .ODT_EN_0                  ( GND_net ), // tied to 1'b0 from definition
        // Outputs
        .TX_0                      ( LANE_2_IOD_DQSW_TRAINING_TX_0 ),
        .OE_0                      ( LANE_2_IOD_DQSW_TRAINING_OE_0 ),
        .DELAY_LINE_OUT_OF_RANGE_0 ( LANE_2_IOD_DQSW_TRAINING_DELAY_LINE_OUT_OF_RANGE_0 ),
        .EYE_MONITOR_EARLY_0       ( LANE_2_IOD_DQSW_TRAINING_EYE_MONITOR_EARLY_0 ),
        .EYE_MONITOR_LATE_0        ( LANE_2_IOD_DQSW_TRAINING_EYE_MONITOR_LATE_0 ),
        .RX_DATA_0                 ( RX_DATA_0_net_10 ) 
        );

//--------PF_DDR4_SS_DDRPHY_BLK_LANE_2_IOD_READ_TRAINING_PF_IOD   -   Actel:SgCore:PF_IOD:1.0.218
PF_DDR4_SS_DDRPHY_BLK_LANE_2_IOD_READ_TRAINING_PF_IOD LANE_2_IOD_READ_TRAINING(
        // Inputs
        .RX_P_0                    ( LANE_2_IOD_DQS_DQS_N ),
        .ARST_N                    ( LANE_2_CTRL_ARST_N ),
        .RX_SYNC_RST               ( LANE_2_CTRL_RX_SYNC_RST ),
        .TX_SYNC_RST               ( LANE_2_CTRL_TX_SYNC_RST ),
        .HS_IO_CLK                 ( HS_IO_CLK ),
        .TX_DQS                    ( LANE_2_CTRL_TX_DQS ),
        .FIFO_WR_PTR               ( LANE_2_CTRL_FIFO_WR_PTR ),
        .FIFO_RD_PTR               ( LANE_2_CTRL_FIFO_RD_PTR ),
        .TX_DATA_0                 ( TX_DATA_0_net_21 ),
        .OE_DATA_0                 ( OE_DATA_0_net_12 ),
        .EYE_MONITOR_CLEAR_FLAGS_0 ( IOD_TRAINING_0_DQSW270_EYE_MONITOR_CLR_FLAGS2to2 ),
        .DELAY_LINE_MOVE_0         ( IOD_TRAINING_0_DQSW270_DELAY_LINE_MOVE2to2 ),
        .DELAY_LINE_DIRECTION_0    ( IOD_TRAINING_0_DQSW270_DELAY_LINE_DIRECTION2to2 ),
        .DELAY_LINE_LOAD_0         ( IOD_TRAINING_0_DQSW270_DELAY_LINE_LOAD2to2 ),
        .FAB_CLK                   ( SYS_CLK ),
        .ODT_EN_0                  ( GND_net ), // tied to 1'b0 from definition
        // Outputs
        .DELAY_LINE_OUT_OF_RANGE_0 ( LANE_2_IOD_READ_TRAINING_DELAY_LINE_OUT_OF_RANGE_0 ),
        .EYE_MONITOR_EARLY_0       ( LANE_2_IOD_READ_TRAINING_EYE_MONITOR_EARLY_0 ),
        .EYE_MONITOR_LATE_0        ( LANE_2_IOD_READ_TRAINING_EYE_MONITOR_LATE_0 ),
        .RX_DATA_0                 ( RX_DATA_0_net_11 ),
        .DDR_DO_READ               ( LANE_2_IOD_READ_TRAINING_DDR_DO_READ ),
        .SWITCH                    ( LANE_2_IOD_READ_TRAINING_SWITCH ) 
        );

//--------PF_DDR4_SS_DDRPHY_BLK_LANE_3_CTRL_PF_LANECTRL   -   Actel:SgCore:PF_LANECTRL:2.0.102
PF_DDR4_SS_DDRPHY_BLK_LANE_3_CTRL_PF_LANECTRL LANE_3_CTRL(
        // Inputs
        .DQS                        ( LANE_3_IOD_DQS_DQS ),
        .HS_IO_CLK                  ( HS_IO_CLK_net_3 ),
        .DLL_CODE                   ( DLL_CODE ),
        .FAB_CLK                    ( SYS_CLK ),
        .RESET                      ( SYNC_SYS_RST_N_net_0 ),
        .DDR_READ                   ( DFI_RDLVL_GATE_EN ),
        .READ_CLK_SEL               ( READ_CLK_SEL_net_3 ),
        .DELAY_LINE_SEL             ( IOD_TRAINING_0_DELAY_LINE_SEL_RD3to3 ),
        .DELAY_LINE_LOAD            ( IOD_TRAINING_0_LOAD35to35 ),
        .DELAY_LINE_DIRECTION       ( IOD_TRAINING_0_DIRECTION35to35 ),
        .DELAY_LINE_MOVE            ( IOD_TRAINING_0_MOVE35to35 ),
        .HS_IO_CLK_PAUSE            ( IOD_TRAINING_0_INIT_PAUSE3to3 ),
        .EYE_MONITOR_WIDTH_IN       ( EYE_MONITOR_WIDTH_IN_const_net_3 ),
        .ODT_EN                     ( VCC_net ),
        .CDR_CLK_A_SEL              ( IOD_TRAINING_0_DQSW_SELA31to24 ),
        .DDR_DO_READ                ( LANE_3_IOD_READ_TRAINING_DDR_DO_READ ),
        .SWITCH                     ( LANE_3_IOD_READ_TRAINING_SWITCH ),
        // Outputs
        .EYE_MONITOR_WIDTH_OUT      ( LANE_3_CTRL_EYE_MONITOR_WIDTH_OUT ),
        .ODT_EN_SEL                 (  ),
        .RX_DQS_90                  ( LANE_3_CTRL_RX_DQS_90 ),
        .TX_DQS                     ( LANE_3_CTRL_TX_DQS ),
        .TX_DQS_270                 ( LANE_3_CTRL_TX_DQS_270 ),
        .FIFO_WR_PTR                ( LANE_3_CTRL_FIFO_WR_PTR ),
        .FIFO_RD_PTR                ( LANE_3_CTRL_FIFO_RD_PTR ),
        .ARST_N                     ( LANE_3_CTRL_ARST_N ),
        .RX_SYNC_RST                ( LANE_3_CTRL_RX_SYNC_RST ),
        .TX_SYNC_RST                ( LANE_3_CTRL_TX_SYNC_RST ),
        .ODT_EN_OUT                 (  ),
        .RX_DATA_VALID              ( LANE_3_CTRL_RX_DATA_VALID ),
        .RX_BURST_DETECT            ( LANE_3_CTRL_RX_BURST_DETECT ),
        .RX_DELAY_LINE_OUT_OF_RANGE ( LANE_3_CTRL_RX_DELAY_LINE_OUT_OF_RANGE ),
        .TX_DELAY_LINE_OUT_OF_RANGE ( LANE_3_CTRL_TX_DELAY_LINE_OUT_OF_RANGE ),
        .A_OUT_RST_N                (  ) 
        );

//--------PF_DDR4_SS_DDRPHY_BLK_LANE_3_IOD_DM_PF_IOD   -   Actel:SgCore:PF_IOD:1.0.218
PF_DDR4_SS_DDRPHY_BLK_LANE_3_IOD_DM_PF_IOD LANE_3_IOD_DM(
        // Inputs
        .ARST_N                    ( LANE_3_CTRL_ARST_N ),
        .RX_SYNC_RST               ( LANE_3_CTRL_RX_SYNC_RST ),
        .TX_SYNC_RST               ( LANE_3_CTRL_TX_SYNC_RST ),
        .HS_IO_CLK                 ( HS_IO_CLK ),
        .TX_DQS                    ( LANE_3_CTRL_TX_DQS ),
        .TX_DATA_0                 ( TX_DATA_0_net_22 ),
        .OE_DATA_0                 ( OE_DATA_0_net_13 ),
        .DELAY_LINE_MOVE_0         ( GND_net ),
        .DELAY_LINE_DIRECTION_0    ( GND_net ),
        .DELAY_LINE_LOAD_0         ( GND_net ),
        .FAB_CLK                   ( SYS_CLK ),
        .ODT_EN_0                  ( GND_net ), // tied to 1'b0 from definition
        // Outputs
        .DELAY_LINE_OUT_OF_RANGE_0 (  ),
        .PAD_O                     ( DM_N_2 ),
        .RX_FB                     ( LANE_3_IOD_DM_RX_FB ) 
        );

//--------PF_DDR4_SS_DDRPHY_BLK_LANE_3_IOD_DQ_PF_IOD   -   Actel:SgCore:PF_IOD:1.0.218
PF_DDR4_SS_DDRPHY_BLK_LANE_3_IOD_DQ_PF_IOD LANE_3_IOD_DQ(
        // Inputs
        .ARST_N                    ( LANE_3_CTRL_ARST_N ),
        .RX_SYNC_RST               ( LANE_3_CTRL_RX_SYNC_RST ),
        .TX_SYNC_RST               ( LANE_3_CTRL_TX_SYNC_RST ),
        .HS_IO_CLK                 ( HS_IO_CLK ),
        .RX_DQS_90                 ( LANE_3_CTRL_RX_DQS_90 ),
        .TX_DQS                    ( LANE_3_CTRL_TX_DQS ),
        .FIFO_WR_PTR               ( LANE_3_CTRL_FIFO_WR_PTR ),
        .FIFO_RD_PTR               ( LANE_3_CTRL_FIFO_RD_PTR ),
        .EYE_MONITOR_LANE_WIDTH    ( LANE_3_CTRL_EYE_MONITOR_WIDTH_OUT ),
        .TX_DATA_0                 ( TX_DATA_0_net_23 ),
        .TX_DATA_1                 ( TX_DATA_1_net_6 ),
        .TX_DATA_2                 ( TX_DATA_2_net_4 ),
        .TX_DATA_3                 ( TX_DATA_3_net_4 ),
        .TX_DATA_4                 ( TX_DATA_4_net_4 ),
        .TX_DATA_5                 ( TX_DATA_5_net_4 ),
        .TX_DATA_6                 ( TX_DATA_6_net_4 ),
        .TX_DATA_7                 ( TX_DATA_7_net_4 ),
        .OE_DATA_0                 ( OE_DATA_0_net_14 ),
        .OE_DATA_1                 ( OE_DATA_1_net_3 ),
        .OE_DATA_2                 ( OE_DATA_2_net_3 ),
        .OE_DATA_3                 ( OE_DATA_3_net_3 ),
        .OE_DATA_4                 ( OE_DATA_4_net_3 ),
        .OE_DATA_5                 ( OE_DATA_5_net_3 ),
        .OE_DATA_6                 ( OE_DATA_6_net_3 ),
        .OE_DATA_7                 ( OE_DATA_7_net_3 ),
        .EYE_MONITOR_CLEAR_FLAGS_0 ( GND_net ),
        .EYE_MONITOR_CLEAR_FLAGS_1 ( GND_net ),
        .EYE_MONITOR_CLEAR_FLAGS_2 ( GND_net ),
        .EYE_MONITOR_CLEAR_FLAGS_3 ( GND_net ),
        .EYE_MONITOR_CLEAR_FLAGS_4 ( GND_net ),
        .EYE_MONITOR_CLEAR_FLAGS_5 ( GND_net ),
        .EYE_MONITOR_CLEAR_FLAGS_6 ( GND_net ),
        .EYE_MONITOR_CLEAR_FLAGS_7 ( GND_net ),
        .DELAY_LINE_MOVE_0         ( IOD_TRAINING_0_MOVE27to27 ),
        .DELAY_LINE_MOVE_1         ( IOD_TRAINING_0_MOVE28to28 ),
        .DELAY_LINE_MOVE_2         ( IOD_TRAINING_0_MOVE29to29 ),
        .DELAY_LINE_MOVE_3         ( IOD_TRAINING_0_MOVE30to30 ),
        .DELAY_LINE_MOVE_4         ( IOD_TRAINING_0_MOVE31to31 ),
        .DELAY_LINE_MOVE_5         ( IOD_TRAINING_0_MOVE32to32 ),
        .DELAY_LINE_MOVE_6         ( IOD_TRAINING_0_MOVE33to33 ),
        .DELAY_LINE_MOVE_7         ( IOD_TRAINING_0_MOVE34to34 ),
        .DELAY_LINE_DIRECTION_0    ( IOD_TRAINING_0_DIRECTION27to27 ),
        .DELAY_LINE_DIRECTION_1    ( IOD_TRAINING_0_DIRECTION28to28 ),
        .DELAY_LINE_DIRECTION_2    ( IOD_TRAINING_0_DIRECTION29to29 ),
        .DELAY_LINE_DIRECTION_3    ( IOD_TRAINING_0_DIRECTION30to30 ),
        .DELAY_LINE_DIRECTION_4    ( IOD_TRAINING_0_DIRECTION31to31 ),
        .DELAY_LINE_DIRECTION_5    ( IOD_TRAINING_0_DIRECTION32to32 ),
        .DELAY_LINE_DIRECTION_6    ( IOD_TRAINING_0_DIRECTION33to33 ),
        .DELAY_LINE_DIRECTION_7    ( IOD_TRAINING_0_DIRECTION34to34 ),
        .DELAY_LINE_LOAD_0         ( IOD_TRAINING_0_LOAD27to27 ),
        .DELAY_LINE_LOAD_1         ( IOD_TRAINING_0_LOAD28to28 ),
        .DELAY_LINE_LOAD_2         ( IOD_TRAINING_0_LOAD29to29 ),
        .DELAY_LINE_LOAD_3         ( IOD_TRAINING_0_LOAD30to30 ),
        .DELAY_LINE_LOAD_4         ( IOD_TRAINING_0_LOAD31to31 ),
        .DELAY_LINE_LOAD_5         ( IOD_TRAINING_0_LOAD32to32 ),
        .DELAY_LINE_LOAD_6         ( IOD_TRAINING_0_LOAD33to33 ),
        .DELAY_LINE_LOAD_7         ( IOD_TRAINING_0_LOAD34to34 ),
        .FAB_CLK                   ( SYS_CLK ),
        .ODT_EN_0                  ( GND_net ), // tied to 1'b0 from definition
        .ODT_EN_1                  ( GND_net ), // tied to 1'b0 from definition
        .ODT_EN_2                  ( GND_net ), // tied to 1'b0 from definition
        .ODT_EN_3                  ( GND_net ), // tied to 1'b0 from definition
        .ODT_EN_4                  ( GND_net ), // tied to 1'b0 from definition
        .ODT_EN_5                  ( GND_net ), // tied to 1'b0 from definition
        .ODT_EN_6                  ( GND_net ), // tied to 1'b0 from definition
        .ODT_EN_7                  ( GND_net ), // tied to 1'b0 from definition
        // Outputs
        .DELAY_LINE_OUT_OF_RANGE_0 ( LANE_3_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_0 ),
        .DELAY_LINE_OUT_OF_RANGE_1 ( LANE_3_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_1 ),
        .DELAY_LINE_OUT_OF_RANGE_2 ( LANE_3_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_2 ),
        .DELAY_LINE_OUT_OF_RANGE_3 ( LANE_3_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_3 ),
        .DELAY_LINE_OUT_OF_RANGE_4 ( LANE_3_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_4 ),
        .DELAY_LINE_OUT_OF_RANGE_5 ( LANE_3_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_5 ),
        .DELAY_LINE_OUT_OF_RANGE_6 ( LANE_3_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_6 ),
        .DELAY_LINE_OUT_OF_RANGE_7 ( LANE_3_IOD_DQ_DELAY_LINE_OUT_OF_RANGE_7 ),
        .EYE_MONITOR_EARLY_0       (  ),
        .EYE_MONITOR_EARLY_1       (  ),
        .EYE_MONITOR_EARLY_2       (  ),
        .EYE_MONITOR_EARLY_3       (  ),
        .EYE_MONITOR_EARLY_4       (  ),
        .EYE_MONITOR_EARLY_5       (  ),
        .EYE_MONITOR_EARLY_6       (  ),
        .EYE_MONITOR_EARLY_7       (  ),
        .EYE_MONITOR_LATE_0        (  ),
        .EYE_MONITOR_LATE_1        (  ),
        .EYE_MONITOR_LATE_2        (  ),
        .EYE_MONITOR_LATE_3        (  ),
        .EYE_MONITOR_LATE_4        (  ),
        .EYE_MONITOR_LATE_5        (  ),
        .EYE_MONITOR_LATE_6        (  ),
        .EYE_MONITOR_LATE_7        (  ),
        .RX_DATA_0                 ( RX_DATA_0_net_12 ),
        .RX_DATA_1                 ( RX_DATA_1_net_3 ),
        .RX_DATA_2                 ( RX_DATA_2_net_3 ),
        .RX_DATA_3                 ( RX_DATA_3_net_3 ),
        .RX_DATA_4                 ( RX_DATA_4_net_3 ),
        .RX_DATA_5                 ( RX_DATA_5_net_3 ),
        .RX_DATA_6                 ( RX_DATA_6_net_3 ),
        .RX_DATA_7                 ( RX_DATA_7_net_3 ),
        .RX_BYPASS_DATA_0          ( LANE_3_IOD_DQ_RX_BYPASS_DATA_0 ),
        .RX_BYPASS_DATA_1          ( LANE_3_IOD_DQ_RX_BYPASS_DATA_1 ),
        .RX_BYPASS_DATA_2          ( LANE_3_IOD_DQ_RX_BYPASS_DATA_2 ),
        .RX_BYPASS_DATA_3          ( LANE_3_IOD_DQ_RX_BYPASS_DATA_3 ),
        .RX_BYPASS_DATA_4          ( LANE_3_IOD_DQ_RX_BYPASS_DATA_4 ),
        .RX_BYPASS_DATA_5          ( LANE_3_IOD_DQ_RX_BYPASS_DATA_5 ),
        .RX_BYPASS_DATA_6          ( LANE_3_IOD_DQ_RX_BYPASS_DATA_6 ),
        .RX_BYPASS_DATA_7          ( LANE_3_IOD_DQ_RX_BYPASS_DATA_7 ),
        // Inouts
        .PAD                       ( { DQ[31:31] , DQ[30:30] , DQ[29:29] , DQ[28:28] , DQ[27:27] , DQ[26:26] , DQ[25:25] , DQ[24:24] } ) 
        );

//--------PF_DDR4_SS_DDRPHY_BLK_LANE_3_IOD_DQS_PF_IOD   -   Actel:SgCore:PF_IOD:1.0.218
PF_DDR4_SS_DDRPHY_BLK_LANE_3_IOD_DQS_PF_IOD LANE_3_IOD_DQS(
        // Inputs
        .ARST_N                    ( LANE_3_CTRL_ARST_N ),
        .RX_SYNC_RST               ( LANE_3_CTRL_RX_SYNC_RST ),
        .TX_SYNC_RST               ( LANE_3_CTRL_TX_SYNC_RST ),
        .HS_IO_CLK                 ( HS_IO_CLK ),
        .RX_DQS_90                 ( LANE_3_CTRL_RX_DQS_90 ),
        .TX_DQS_270                ( LANE_3_CTRL_TX_DQS_270 ),
        .FIFO_WR_PTR               ( LANE_3_CTRL_FIFO_WR_PTR ),
        .FIFO_RD_PTR               ( LANE_3_CTRL_FIFO_RD_PTR ),
        .EYE_MONITOR_LANE_WIDTH    ( LANE_3_CTRL_EYE_MONITOR_WIDTH_OUT ),
        .TX_DATA_0                 ( TX_DATA_0_const_net_6 ),
        .OE_DATA_0                 ( OE_DATA_0_net_15 ),
        .EYE_MONITOR_CLEAR_FLAGS_0 ( GND_net ),
        .DELAY_LINE_MOVE_0         ( GND_net ),
        .DELAY_LINE_DIRECTION_0    ( GND_net ),
        .DELAY_LINE_LOAD_0         ( GND_net ),
        .FAB_CLK                   ( SYS_CLK ),
        .ODT_EN_0                  ( GND_net ), // tied to 1'b0 from definition
        // Outputs
        .DELAY_LINE_OUT_OF_RANGE_0 (  ),
        .EYE_MONITOR_EARLY_0       (  ),
        .EYE_MONITOR_LATE_0        (  ),
        .RX_DATA_0                 (  ),
        .DQS                       ( LANE_3_IOD_DQS_DQS ),
        .DQS_N                     ( LANE_3_IOD_DQS_DQS_N ),
        // Inouts
        .PAD                       ( DQS[3:3] ),
        .PAD_N                     ( DQS_N[3:3] ) 
        );

//--------PF_DDR4_SS_DDRPHY_BLK_LANE_3_IOD_DQSW_TRAINING_PF_IOD   -   Actel:SgCore:PF_IOD:1.0.218
PF_DDR4_SS_DDRPHY_BLK_LANE_3_IOD_DQSW_TRAINING_PF_IOD LANE_3_IOD_DQSW_TRAINING(
        // Inputs
        .RX_N_0                    ( LANE_3_IOD_DM_RX_FB ),
        .HS_IO_CLK                 ( HS_IO_CLK ),
        .TX_DATA_0                 ( TX_DATA_0_const_net_7 ),
        .OE_DATA_0                 ( OE_DATA_0_const_net_15 ),
        .EYE_MONITOR_CLEAR_FLAGS_0 ( IOD_TRAINING_0_DQSW_EYE_MONITOR_CLR_FLAGS3to3 ),
        .DELAY_LINE_MOVE_0         ( IOD_TRAINING_0_DQSW_DELAY_LINE_MOVE3to3 ),
        .DELAY_LINE_DIRECTION_0    ( IOD_TRAINING_0_DQSW_DELAY_LINE_DIRECTION3to3 ),
        .DELAY_LINE_LOAD_0         ( IOD_TRAINING_0_DQSW_DELAY_LINE_LOAD3to3 ),
        .FAB_CLK                   ( SYS_CLK ),
        .ODT_EN_0                  ( GND_net ), // tied to 1'b0 from definition
        // Outputs
        .TX_0                      ( LANE_3_IOD_DQSW_TRAINING_TX_0 ),
        .OE_0                      ( LANE_3_IOD_DQSW_TRAINING_OE_0 ),
        .DELAY_LINE_OUT_OF_RANGE_0 ( LANE_3_IOD_DQSW_TRAINING_DELAY_LINE_OUT_OF_RANGE_0 ),
        .EYE_MONITOR_EARLY_0       ( LANE_3_IOD_DQSW_TRAINING_EYE_MONITOR_EARLY_0 ),
        .EYE_MONITOR_LATE_0        ( LANE_3_IOD_DQSW_TRAINING_EYE_MONITOR_LATE_0 ),
        .RX_DATA_0                 ( RX_DATA_0_net_13 ) 
        );

//--------PF_DDR4_SS_DDRPHY_BLK_LANE_3_IOD_READ_TRAINING_PF_IOD   -   Actel:SgCore:PF_IOD:1.0.218
PF_DDR4_SS_DDRPHY_BLK_LANE_3_IOD_READ_TRAINING_PF_IOD LANE_3_IOD_READ_TRAINING(
        // Inputs
        .RX_P_0                    ( LANE_3_IOD_DQS_DQS_N ),
        .ARST_N                    ( LANE_3_CTRL_ARST_N ),
        .RX_SYNC_RST               ( LANE_3_CTRL_RX_SYNC_RST ),
        .TX_SYNC_RST               ( LANE_3_CTRL_TX_SYNC_RST ),
        .HS_IO_CLK                 ( HS_IO_CLK ),
        .TX_DQS                    ( LANE_3_CTRL_TX_DQS ),
        .FIFO_WR_PTR               ( LANE_3_CTRL_FIFO_WR_PTR ),
        .FIFO_RD_PTR               ( LANE_3_CTRL_FIFO_RD_PTR ),
        .TX_DATA_0                 ( TX_DATA_0_net_24 ),
        .OE_DATA_0                 ( OE_DATA_0_net_16 ),
        .EYE_MONITOR_CLEAR_FLAGS_0 ( IOD_TRAINING_0_DQSW270_EYE_MONITOR_CLR_FLAGS3to3 ),
        .DELAY_LINE_MOVE_0         ( IOD_TRAINING_0_DQSW270_DELAY_LINE_MOVE3to3 ),
        .DELAY_LINE_DIRECTION_0    ( IOD_TRAINING_0_DQSW270_DELAY_LINE_DIRECTION3to3 ),
        .DELAY_LINE_LOAD_0         ( IOD_TRAINING_0_DQSW270_DELAY_LINE_LOAD3to3 ),
        .FAB_CLK                   ( SYS_CLK ),
        .ODT_EN_0                  ( GND_net ), // tied to 1'b0 from definition
        // Outputs
        .DELAY_LINE_OUT_OF_RANGE_0 ( LANE_3_IOD_READ_TRAINING_DELAY_LINE_OUT_OF_RANGE_0 ),
        .EYE_MONITOR_EARLY_0       ( LANE_3_IOD_READ_TRAINING_EYE_MONITOR_EARLY_0 ),
        .EYE_MONITOR_LATE_0        ( LANE_3_IOD_READ_TRAINING_EYE_MONITOR_LATE_0 ),
        .RX_DATA_0                 ( RX_DATA_0_net_14 ),
        .DDR_DO_READ               ( LANE_3_IOD_READ_TRAINING_DDR_DO_READ ),
        .SWITCH                    ( LANE_3_IOD_READ_TRAINING_SWITCH ) 
        );

//--------PF_DDR4_SS_DDRPHY_BLK_LANECTRL_ADDR_CMD_0_PF_LANECTRL   -   Actel:SgCore:PF_LANECTRL:2.0.102
PF_DDR4_SS_DDRPHY_BLK_LANECTRL_ADDR_CMD_0_PF_LANECTRL LANECTRL_ADDR_CMD_0(
        // Inputs
        .HS_IO_CLK                  ( HS_IO_CLK ),
        .DLL_CODE                   ( DLL_CODE ),
        .FAB_CLK                    ( SYS_CLK ),
        .RESET                      ( GND_net ),
        .DDR_READ                   ( GND_net ), // tied to 1'b0 from definition
        .DELAY_LINE_SEL             ( GND_net ), // tied to 1'b0 from definition
        .DELAY_LINE_LOAD            ( VCC_net ),
        .DELAY_LINE_DIRECTION       ( GND_net ), // tied to 1'b0 from definition
        .DELAY_LINE_MOVE            ( GND_net ), // tied to 1'b0 from definition
        .HS_IO_CLK_PAUSE            ( CLKINT_CMD_Y ),
        .EYE_MONITOR_WIDTH_IN       ( EYE_MONITOR_WIDTH_IN_const_net_4 ), // tied to 3'h0 from definition
        .CDR_CLK_A_SEL              ( CDR_CLK_A_SEL_const_net_0 ), // tied to 8'h00 from definition
        // Outputs
        .EYE_MONITOR_WIDTH_OUT      (  ),
        .RX_DQS_90                  (  ),
        .TX_DQS                     (  ),
        .TX_DQS_270                 ( LANECTRL_ADDR_CMD_0_TX_DQS_270 ),
        .FIFO_WR_PTR                (  ),
        .FIFO_RD_PTR                (  ),
        .ARST_N                     ( LANECTRL_ADDR_CMD_0_ARST_N ),
        .RX_SYNC_RST                ( LANECTRL_ADDR_CMD_0_RX_SYNC_RST ),
        .TX_SYNC_RST                ( LANECTRL_ADDR_CMD_0_TX_SYNC_RST ),
        .RX_DATA_VALID              (  ),
        .RX_BURST_DETECT            (  ),
        .RX_DELAY_LINE_OUT_OF_RANGE (  ),
        .TX_DELAY_LINE_OUT_OF_RANGE (  ),
        .A_OUT_RST_N                (  ) 
        );

//--------OUTBUF_FEEDBACK
OUTBUF_FEEDBACK OB_A_12(
        // Inputs
        .D   ( IOD_A_12_TX_0 ),
        // Outputs
        .Y   ( OB_A_12_Y ),
        .PAD ( A_11 ) 
        );

//--------OUTBUF_FEEDBACK_DIFF
OUTBUF_FEEDBACK_DIFF OB_DIFF_CK0(
        // Inputs
        .D    ( REF_CLK ),
        // Outputs
        .Y    ( OB_DIFF_CK0_Y ),
        .PADP ( CK0_net_0 ),
        .PADN ( CK0_N_net_0 ) 
        );

//--------TRIBUFF
TRIBUFF TRI_SHIELD_0(
        // Inputs
        .D   ( LANE_0_IOD_DQSW_TRAINING_TX_0 ),
        .E   ( LANE_0_IOD_DQSW_TRAINING_OE_0 ),
        // Outputs
        .PAD ( SHIELD0_net_0 ) 
        );

//--------TRIBUFF
TRIBUFF TRI_SHIELD_1(
        // Inputs
        .D   ( LANE_1_IOD_DQSW_TRAINING_TX_0 ),
        .E   ( LANE_1_IOD_DQSW_TRAINING_OE_0 ),
        // Outputs
        .PAD ( SHIELD1_net_0 ) 
        );

//--------TRIBUFF
TRIBUFF TRI_SHIELD_2(
        // Inputs
        .D   ( LANE_2_IOD_DQSW_TRAINING_TX_0 ),
        .E   ( LANE_2_IOD_DQSW_TRAINING_OE_0 ),
        // Outputs
        .PAD ( SHIELD2_net_0 ) 
        );

//--------TRIBUFF
TRIBUFF TRI_SHIELD_3(
        // Inputs
        .D   ( LANE_3_IOD_DQSW_TRAINING_TX_0 ),
        .E   ( LANE_3_IOD_DQSW_TRAINING_OE_0 ),
        // Outputs
        .PAD ( SHIELD3_net_0 ) 
        );


endmodule
