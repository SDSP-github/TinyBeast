`timescale 1ns/1ps
// ****************************************************************************/
// Microsemi Corporation Proprietary and Confidential
// Copyright 2017 Microsemi Corporation.  All rights reserved.
//
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
// ACCORDANCE WITH THE MICROSEMI LICENSE AGREEMENT AND MUST BE APPROVED
// IN ADVANCE IN WRITING.
//
// Description: 
//
// SVN Revision Information:
// SVN $Revision: 37592 $
// SVN $Date: 2021-02-02 23:05:01 +0530 (Tue, 02 Feb 2021) $
//
// Resolved SARs
// SAR      Date     Who   Description
//
// Notes:
//
// ****************************************************************************/
//`define TEST_CASE_0 1
//`define TEST_CASE_1 1
module AXI4StreamMaster (
    // General inputs
    clock,
    resetn,
    
    // AXI4Stream inputs
    TREADY,
    
    // AXI4Stream outputs
    TVALID,
    TID,
    TSTRB,
    TKEEP,
    TLAST,
    TDATA,
    TDEST
);

////////////////////////////////////////////////////////////////////////////////
// Parameters
////////////////////////////////////////////////////////////////////////////////
parameter ADDR_WIDTH    = 10;
parameter DATA_WIDTH    = 32;
parameter RAM_INIT_FILE = "./ram_init.mem";
parameter ID_WIDTH      = 2;

////////////////////////////////////////////////////////////////////////////////
// Port directions
////////////////////////////////////////////////////////////////////////////////
// General inputs
input                               clock;
input                               resetn;
    
// AXI4Stream inputs
input                               TREADY;

// AXI4Stream outputs
output reg                          TVALID;
output reg                          TID;
output reg  [(DATA_WIDTH/8)-1:0]    TSTRB;
output reg  [(DATA_WIDTH/8)-1:0]    TKEEP;
output reg                          TLAST;
output reg  [DATA_WIDTH-1:0]        TDATA;
output reg  [1:0]                   TDEST;

////////////////////////////////////////////////////////////////////////////////
// Internal signals
////////////////////////////////////////////////////////////////////////////////
reg  [ADDR_WIDTH-1:0]               rdAddr;
wire [DATA_WIDTH-1:0]               rdData;
reg  [7:0]                          RAM_BUFFER [0:(2**ADDR_WIDTH)-1];

// Initialize the stream interface outputs
initial
    begin
        TVALID = 1'b0;
        TLAST  = 1'b0;
        TID    = {ID_WIDTH{1'b0}};
        TDATA  = {DATA_WIDTH{1'b0}};
        TSTRB  = {(DATA_WIDTH/8){1'b0}};
        TKEEP  = {(DATA_WIDTH/8){1'b0}};
        TDEST  = 2'b0;
    end

// Initialize the contents of the RAM for simulation
initial
    begin
        $readmemb(RAM_INIT_FILE, RAM_BUFFER); 
    end
    
////////////////////////////////////////////////////////////////////////////////
// Asynchronous read
////////////////////////////////////////////////////////////////////////////////
generate
    genvar  read_offset;
    for(read_offset=0; read_offset<(DATA_WIDTH/8); read_offset = read_offset + 1)
        begin : mem_read
            assign rdData[(((read_offset+1)<<3)-1):(read_offset<<3)] = RAM_BUFFER[(rdAddr+read_offset)]; 
        end
endgenerate

////////////////////////////////////////////////////////////////////////////////
// Stream write task
////////////////////////////////////////////////////////////////////////////////
task axi4_stream_write;
    input [1:0]                         destRouteInfo;
    input [23:0]                        dstNumOfBytes;
    input [31:0]                        srcAddr;
    integer                             offset;
    integer                             byteCnt;
    integer                             trigger;
    integer                             cycleCnt;
    begin
        // Initialize variables
        offset  = 0;
        byteCnt = 0;
        rdAddr  = 0;
        cycleCnt = 0;
        // Wait for a clock edge before we start driving out data
        @(posedge clock);
        if (dstNumOfBytes > (DATA_WIDTH/8))
            begin
                // More than 4 bytes in the entire stream transaction
                while((dstNumOfBytes - byteCnt) > (DATA_WIDTH/8))
                    begin
                        // More than one transfer in the stream transaction
                        // This is not the first or the last transfer so all byte
                        // lanes contain valid data
                        offset  = offset + (DATA_WIDTH/8);
                        TVALID  = 1'b1;
                        TLAST   = 1'b0;
                        TID     = {ID_WIDTH{1'b0}};
                        TDATA   = rdData;
                        TSTRB   = {(DATA_WIDTH/8){1'b1}};
                        TKEEP   = {(DATA_WIDTH/8){1'b1}};
                        TDEST   = destRouteInfo;
                        byteCnt = byteCnt + (DATA_WIDTH/8);
                        trigger = 0;
                        while (trigger != 1) begin
                            @ (posedge clock);
                            trigger = TREADY;
                        end
                        cycleCnt = cycleCnt + 1;
                        rdAddr  = srcAddr + offset;
                        #1;
                    end
            end
        // Last beat coming out or transfer consists of a single beat
        TVALID = 1'b1;
        TLAST  = 1'b1;
        TID    = {ID_WIDTH{1'b0}};
        TDATA  = rdData;
        if (DATA_WIDTH == 32)
            begin
                TSTRB  = ((dstNumOfBytes[1:0]) == 1) ? 4'b0001 :
                         ((dstNumOfBytes[1:0]) == 2) ? 4'b0011 :
                         ((dstNumOfBytes[1:0]) == 3) ? 4'b0111 :
                         4'b1111;
            end
        else if (DATA_WIDTH == 64)
            begin
                TSTRB = ((dstNumOfBytes[2:0]) == 1) ? 8'b0000_0001 :
                        ((dstNumOfBytes[2:0]) == 2) ? 8'b0000_0011 :
                        ((dstNumOfBytes[2:0]) == 3) ? 8'b0000_0111 :
                        ((dstNumOfBytes[2:0]) == 4) ? 8'b0000_1111 :
                        ((dstNumOfBytes[2:0]) == 5) ? 8'b0001_1111 :
                        ((dstNumOfBytes[2:0]) == 6) ? 8'b0011_1111 :
                        ((dstNumOfBytes[2:0]) == 7) ? 8'b0111_1111 :
                        8'b1111_1111;
            end
        else if (DATA_WIDTH == 128)
            begin
                TSTRB = ((dstNumOfBytes[3:0]) == 1)  ? 16'b0000_0000_0000_0001 :
                        ((dstNumOfBytes[3:0]) == 2)  ? 16'b0000_0000_0000_0011 :
                        ((dstNumOfBytes[3:0]) == 3)  ? 16'b0000_0000_0000_0111 :
                        ((dstNumOfBytes[3:0]) == 4)  ? 16'b0000_0000_0000_1111 :
                        ((dstNumOfBytes[3:0]) == 5)  ? 16'b0000_0000_0001_1111 :
                        ((dstNumOfBytes[3:0]) == 6)  ? 16'b0000_0000_0011_1111 :
                        ((dstNumOfBytes[3:0]) == 7)  ? 16'b0000_0000_0111_1111 :
                        ((dstNumOfBytes[3:0]) == 8)  ? 16'b0000_0000_1111_1111 :
                        ((dstNumOfBytes[3:0]) == 9)  ? 16'b0000_0001_1111_1111 :
                        ((dstNumOfBytes[3:0]) == 10) ? 16'b0000_0011_1111_1111 :
                        ((dstNumOfBytes[3:0]) == 11) ? 16'b0000_0111_1111_1111 :
                        ((dstNumOfBytes[3:0]) == 12) ? 16'b0000_1111_1111_1111 :
                        ((dstNumOfBytes[3:0]) == 13) ? 16'b0001_1111_1111_1111 :
                        ((dstNumOfBytes[3:0]) == 14) ? 16'b0011_1111_1111_1111 :
                        ((dstNumOfBytes[3:0]) == 15) ? 16'b0111_1111_1111_1111 :
                        16'b1111_1111_1111_1111;
            end
        else if (DATA_WIDTH == 256)
            begin
                TSTRB = ((dstNumOfBytes[4:0]) == 1)  ? 32'b0000_0000_0000_0000_0000_0000_0000_0001 :
                        ((dstNumOfBytes[4:0]) == 2)  ? 32'b0000_0000_0000_0000_0000_0000_0000_0011 :
                        ((dstNumOfBytes[4:0]) == 3)  ? 32'b0000_0000_0000_0000_0000_0000_0000_0111 :
                        ((dstNumOfBytes[4:0]) == 4)  ? 32'b0000_0000_0000_0000_0000_0000_0000_1111 :
                        ((dstNumOfBytes[4:0]) == 5)  ? 32'b0000_0000_0000_0000_0000_0000_0001_1111 :
                        ((dstNumOfBytes[4:0]) == 6)  ? 32'b0000_0000_0000_0000_0000_0000_0011_1111 :
                        ((dstNumOfBytes[4:0]) == 7)  ? 32'b0000_0000_0000_0000_0000_0000_0111_1111 :
                        ((dstNumOfBytes[4:0]) == 8)  ? 32'b0000_0000_0000_0000_0000_0000_1111_1111 :
                        ((dstNumOfBytes[4:0]) == 9)  ? 32'b0000_0000_0000_0000_0000_0001_1111_1111 :
                        ((dstNumOfBytes[4:0]) == 10) ? 32'b0000_0000_0000_0000_0000_0011_1111_1111 :
                        ((dstNumOfBytes[4:0]) == 11) ? 32'b0000_0000_0000_0000_0000_0111_1111_1111 :
                        ((dstNumOfBytes[4:0]) == 12) ? 32'b0000_0000_0000_0000_0000_1111_1111_1111 :
                        ((dstNumOfBytes[4:0]) == 13) ? 32'b0000_0000_0000_0000_0001_1111_1111_1111 :
                        ((dstNumOfBytes[4:0]) == 14) ? 32'b0000_0000_0000_0000_0011_1111_1111_1111 :
                        ((dstNumOfBytes[4:0]) == 15) ? 32'b0000_0000_0000_0000_0111_1111_1111_1111 :
                        ((dstNumOfBytes[4:0]) == 16) ? 32'b0000_0000_0000_0000_1111_1111_1111_1111 :
                        ((dstNumOfBytes[4:0]) == 17) ? 32'b0000_0000_0000_0001_1111_1111_1111_1111 :
                        ((dstNumOfBytes[4:0]) == 18) ? 32'b0000_0000_0000_0011_1111_1111_1111_1111 :
                        ((dstNumOfBytes[4:0]) == 19) ? 32'b0000_0000_0000_0111_1111_1111_1111_1111 :
                        ((dstNumOfBytes[4:0]) == 20) ? 32'b0000_0000_0000_1111_1111_1111_1111_1111 :
                        ((dstNumOfBytes[4:0]) == 21) ? 32'b0000_0000_0001_1111_1111_1111_1111_1111 :
                        ((dstNumOfBytes[4:0]) == 22) ? 32'b0000_0000_0011_1111_1111_1111_1111_1111 :
                        ((dstNumOfBytes[4:0]) == 23) ? 32'b0000_0000_0111_1111_1111_1111_1111_1111 :
                        ((dstNumOfBytes[4:0]) == 24) ? 32'b0000_0000_1111_1111_1111_1111_1111_1111 :
                        ((dstNumOfBytes[4:0]) == 25) ? 32'b0000_0001_1111_1111_1111_1111_1111_1111 :
                        ((dstNumOfBytes[4:0]) == 26) ? 32'b0000_0011_1111_1111_1111_1111_1111_1111 :
                        ((dstNumOfBytes[4:0]) == 27) ? 32'b0000_0111_1111_1111_1111_1111_1111_1111 :
                        ((dstNumOfBytes[4:0]) == 28) ? 32'b0000_1111_1111_1111_1111_1111_1111_1111 :
                        ((dstNumOfBytes[4:0]) == 29) ? 32'b0001_1111_1111_1111_1111_1111_1111_1111 :
                        ((dstNumOfBytes[4:0]) == 30) ? 32'b0011_1111_1111_1111_1111_1111_1111_1111 :
                        ((dstNumOfBytes[4:0]) == 31) ? 32'b0111_1111_1111_1111_1111_1111_1111_1111 :
                        32'b1111_1111_1111_1111_1111_1111_1111_1111;
            end
        else if (DATA_WIDTH == 512)
            begin
                TSTRB = ((dstNumOfBytes[5:0]) == 1)  ? 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001 :
                        ((dstNumOfBytes[5:0]) == 2)  ? 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0011 :
                        ((dstNumOfBytes[5:0]) == 3)  ? 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0111 :
                        ((dstNumOfBytes[5:0]) == 4)  ? 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1111 :
                        ((dstNumOfBytes[5:0]) == 5)  ? 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_1111 :
                        ((dstNumOfBytes[5:0]) == 6)  ? 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0011_1111 :
                        ((dstNumOfBytes[5:0]) == 7)  ? 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0111_1111 :
                        ((dstNumOfBytes[5:0]) == 8)  ? 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1111_1111 :
                        ((dstNumOfBytes[5:0]) == 9)  ? 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_1111_1111 :
                        ((dstNumOfBytes[5:0]) == 10) ? 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0011_1111_1111 :
                        ((dstNumOfBytes[5:0]) == 11) ? 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0111_1111_1111 :
                        ((dstNumOfBytes[5:0]) == 12) ? 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1111_1111_1111 :
                        ((dstNumOfBytes[5:0]) == 13) ? 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_1111_1111_1111 :
                        ((dstNumOfBytes[5:0]) == 14) ? 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0011_1111_1111_1111 :
                        ((dstNumOfBytes[5:0]) == 15) ? 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0111_1111_1111_1111 :
                        ((dstNumOfBytes[5:0]) == 16) ? 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1111_1111_1111_1111 :
                        ((dstNumOfBytes[5:0]) == 17) ? 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_1111_1111_1111_1111 :
                        ((dstNumOfBytes[5:0]) == 18) ? 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0011_1111_1111_1111_1111 :
                        ((dstNumOfBytes[5:0]) == 19) ? 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0111_1111_1111_1111_1111 :
                        ((dstNumOfBytes[5:0]) == 20) ? 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1111_1111_1111_1111_1111 :
                        ((dstNumOfBytes[5:0]) == 21) ? 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_1111_1111_1111_1111_1111 :
                        ((dstNumOfBytes[5:0]) == 22) ? 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0011_1111_1111_1111_1111_1111 :
                        ((dstNumOfBytes[5:0]) == 23) ? 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0111_1111_1111_1111_1111_1111 :
                        ((dstNumOfBytes[5:0]) == 24) ? 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1111_1111_1111_1111_1111_1111 :
                        ((dstNumOfBytes[5:0]) == 25) ? 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_1111_1111_1111_1111_1111_1111 :
                        ((dstNumOfBytes[5:0]) == 26) ? 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0011_1111_1111_1111_1111_1111_1111 :
                        ((dstNumOfBytes[5:0]) == 27) ? 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0111_1111_1111_1111_1111_1111_1111 :
                        ((dstNumOfBytes[5:0]) == 28) ? 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_1111_1111_1111_1111_1111_1111_1111 :
                        ((dstNumOfBytes[5:0]) == 29) ? 64'b0000_0000_0000_0000_0000_0000_0000_0000_0001_1111_1111_1111_1111_1111_1111_1111 :
                        ((dstNumOfBytes[5:0]) == 30) ? 64'b0000_0000_0000_0000_0000_0000_0000_0000_0011_1111_1111_1111_1111_1111_1111_1111 :
                        ((dstNumOfBytes[5:0]) == 31) ? 64'b0000_0000_0000_0000_0000_0000_0000_0000_0111_1111_1111_1111_1111_1111_1111_1111 :
                        ((dstNumOfBytes[5:0]) == 32) ? 64'b0000_0000_0000_0000_0000_0000_0000_0000_1111_1111_1111_1111_1111_1111_1111_1111 :
                        ((dstNumOfBytes[5:0]) == 33) ? 64'b0000_0000_0000_0000_0000_0000_0000_0001_1111_1111_1111_1111_1111_1111_1111_1111 :
                        ((dstNumOfBytes[5:0]) == 34) ? 64'b0000_0000_0000_0000_0000_0000_0000_0011_1111_1111_1111_1111_1111_1111_1111_1111 :
                        ((dstNumOfBytes[5:0]) == 35) ? 64'b0000_0000_0000_0000_0000_0000_0000_0111_1111_1111_1111_1111_1111_1111_1111_1111 :
                        ((dstNumOfBytes[5:0]) == 36) ? 64'b0000_0000_0000_0000_0000_0000_0000_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
                        ((dstNumOfBytes[5:0]) == 37) ? 64'b0000_0000_0000_0000_0000_0000_0001_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
                        ((dstNumOfBytes[5:0]) == 38) ? 64'b0000_0000_0000_0000_0000_0000_0011_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
                        ((dstNumOfBytes[5:0]) == 39) ? 64'b0000_0000_0000_0000_0000_0000_0111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
                        ((dstNumOfBytes[5:0]) == 40) ? 64'b0000_0000_0000_0000_0000_0000_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
                        ((dstNumOfBytes[5:0]) == 41) ? 64'b0000_0000_0000_0000_0000_0001_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
                        ((dstNumOfBytes[5:0]) == 42) ? 64'b0000_0000_0000_0000_0000_0011_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
                        ((dstNumOfBytes[5:0]) == 43) ? 64'b0000_0000_0000_0000_0000_0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
                        ((dstNumOfBytes[5:0]) == 44) ? 64'b0000_0000_0000_0000_0000_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
                        ((dstNumOfBytes[5:0]) == 45) ? 64'b0000_0000_0000_0000_0001_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
                        ((dstNumOfBytes[5:0]) == 46) ? 64'b0000_0000_0000_0000_0011_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
                        ((dstNumOfBytes[5:0]) == 47) ? 64'b0000_0000_0000_0000_0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
                        ((dstNumOfBytes[5:0]) == 48) ? 64'b0000_0000_0000_0000_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
                        ((dstNumOfBytes[5:0]) == 49) ? 64'b0000_0000_0000_0001_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
                        ((dstNumOfBytes[5:0]) == 50) ? 64'b0000_0000_0000_0011_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
                        ((dstNumOfBytes[5:0]) == 51) ? 64'b0000_0000_0000_0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
                        ((dstNumOfBytes[5:0]) == 52) ? 64'b0000_0000_0000_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
                        ((dstNumOfBytes[5:0]) == 53) ? 64'b0000_0000_0001_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
                        ((dstNumOfBytes[5:0]) == 54) ? 64'b0000_0000_0011_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
                        ((dstNumOfBytes[5:0]) == 55) ? 64'b0000_0000_0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
                        ((dstNumOfBytes[5:0]) == 56) ? 64'b0000_0000_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
                        ((dstNumOfBytes[5:0]) == 57) ? 64'b0000_0001_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
                        ((dstNumOfBytes[5:0]) == 58) ? 64'b0000_0011_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
                        ((dstNumOfBytes[5:0]) == 59) ? 64'b0000_0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
                        ((dstNumOfBytes[5:0]) == 60) ? 64'b0000_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
                        ((dstNumOfBytes[5:0]) == 61) ? 64'b0001_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
                        ((dstNumOfBytes[5:0]) == 62) ? 64'b0011_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
                        ((dstNumOfBytes[5:0]) == 63) ? 64'b0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111 :
                        64'b1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111;
            end
        TKEEP  = TSTRB;
        TDEST  = destRouteInfo;
        trigger = 0;
        while (trigger != 1) begin
            @ (posedge clock);
            trigger = TREADY;
        end
        // Transaction complete, drive all signals low 
        rdAddr = {ADDR_WIDTH{1'b0}};
        TVALID = 1'b0;
        TLAST  = 1'b0;
        TID    = {ID_WIDTH{1'b0}};
        TDATA  = {DATA_WIDTH{1'b0}};
        TSTRB  = {(DATA_WIDTH/8){1'b0}};
        TKEEP  = {(DATA_WIDTH/8){1'b0}};
        TDEST  = 2'b0;
    end
endtask // axi4_stream_write
    
initial
    begin
        // Wait for the system to come out of reset
        @(posedge resetn);
        #21;
        `include "./axi4_stream_master_application.v"
        $display ($time, "AXI4-Stream write complete");
        // This process doesn't terminate the simulation
    end

endmodule // AXI4StreamMaster