//////////////////////////////////////////////////////////////////////
// Created by SmartDesign Sat Nov  9 06:54:37 2019
// Version: v12.2 12.700.0.21
//////////////////////////////////////////////////////////////////////

`timescale 1ns / 100ps

// tpsram
module tpsram(
    // Inputs
    CLK,
    R_ADDR,
    W_ADDR,
    W_DATA,
    W_EN,
    // Outputs
    R_DATA
);

//--------------------------------------------------------------------
// Input
//--------------------------------------------------------------------
input         CLK;
input  [11:0] R_ADDR;
input  [8:0]  W_ADDR;
input  [63:0] W_DATA;
input         W_EN;
//--------------------------------------------------------------------
// Output
//--------------------------------------------------------------------
output [7:0]  R_DATA;
//--------------------------------------------------------------------
// Nets
//--------------------------------------------------------------------
wire          CLK;
wire   [11:0] R_ADDR;
wire   [7:0]  R_DATA_0;
wire   [8:0]  W_ADDR;
wire   [63:0] W_DATA;
wire          W_EN;
wire   [7:0]  R_DATA_0_net_0;
//--------------------------------------------------------------------
// TiedOff Nets
//--------------------------------------------------------------------
wire          GND_net;
//--------------------------------------------------------------------
// Constant assignments
//--------------------------------------------------------------------
assign GND_net    = 1'b0;
//--------------------------------------------------------------------
// Top level output port assignments
//--------------------------------------------------------------------
assign R_DATA_0_net_0 = R_DATA_0;
assign R_DATA[7:0]    = R_DATA_0_net_0;
//--------------------------------------------------------------------
// Component instances
//--------------------------------------------------------------------
//--------tpsram_tpsram_0_PF_TPSRAM   -   Actel:SgCore:PF_TPSRAM:1.1.108
tpsram_tpsram_0_PF_TPSRAM tpsram_0(
        // Inputs
        .W_DATA ( W_DATA ),
        .W_ADDR ( W_ADDR ),
        .R_ADDR ( R_ADDR ),
        .W_EN   ( W_EN ),
        .CLK    ( CLK ),
        // Outputs
        .R_DATA ( R_DATA_0 ) 
        );


endmodule
