`timescale 1 ns/100 ps
// Version: v2021.2 2021.2.0.11


module PCIe_EP_PCIex4_0_PF_PCIE(
       APB_S_PRDATA,
       APB_S_PREADY,
       APB_S_PSLVERR,
       APB_S_PADDR,
       APB_S_PENABLE,
       APB_S_PSEL,
       APB_S_PWDATA,
       APB_S_PWRITE,
       APB_S_PCLK,
       APB_S_PRESET_N,
       PCIESS_LANE_RXD2_P,
       PCIESS_LANE_RXD2_N,
       PCIESS_LANE_TXD2_P,
       PCIESS_LANE_TXD2_N,
       AXI_CLK,
       AXI_CLK_STABLE,
       PCIE_1_LTSSM,
       PCIE_1_INTERRUPT_OUT,
       PCIE_1_INTERRUPT,
       PCIE_1_TL_CLK_125MHz,
       PCIE_1_M_WDERR,
       PCIE_1_S_RDERR,
       PCIE_1_M_RDERR,
       PCIE_1_S_WDERR,
       PCIE_1_L2_EXIT,
       PCIE_1_HOT_RST_EXIT,
       PCIE_1_DLUP_EXIT,
       PCIE_1_PERST_N,
       PCIESS_AXI_1_M_ARID,
       PCIESS_AXI_1_M_AWID,
       PCIESS_AXI_1_M_ARADDR,
       PCIESS_AXI_1_M_ARBURST,
       PCIESS_AXI_1_M_ARLEN,
       PCIESS_AXI_1_M_ARSIZE,
       PCIESS_AXI_1_M_ARVALID,
       PCIESS_AXI_1_M_AWADDR,
       PCIESS_AXI_1_M_AWBURST,
       PCIESS_AXI_1_M_AWLEN,
       PCIESS_AXI_1_M_AWSIZE,
       PCIESS_AXI_1_M_AWVALID,
       PCIESS_AXI_1_M_BREADY,
       PCIESS_AXI_1_M_RREADY,
       PCIESS_AXI_1_M_WLAST,
       PCIESS_AXI_1_M_WSTRB,
       PCIESS_AXI_1_M_WVALID,
       PCIESS_AXI_1_S_ARREADY,
       PCIESS_AXI_1_S_AWREADY,
       PCIESS_AXI_1_S_BID,
       PCIESS_AXI_1_S_BRESP,
       PCIESS_AXI_1_S_BVALID,
       PCIESS_AXI_1_S_RID,
       PCIESS_AXI_1_S_RLAST,
       PCIESS_AXI_1_S_RRESP,
       PCIESS_AXI_1_S_RVALID,
       PCIESS_AXI_1_S_WREADY,
       PCIESS_AXI_1_M_ARREADY,
       PCIESS_AXI_1_M_AWREADY,
       PCIESS_AXI_1_M_BID,
       PCIESS_AXI_1_M_BRESP,
       PCIESS_AXI_1_M_BVALID,
       PCIESS_AXI_1_M_RID,
       PCIESS_AXI_1_M_RLAST,
       PCIESS_AXI_1_M_RRESP,
       PCIESS_AXI_1_M_RVALID,
       PCIESS_AXI_1_M_WREADY,
       PCIESS_AXI_1_S_ARADDR,
       PCIESS_AXI_1_S_ARBURST,
       PCIESS_AXI_1_S_ARID,
       PCIESS_AXI_1_S_ARLEN,
       PCIESS_AXI_1_S_ARSIZE,
       PCIESS_AXI_1_S_ARVALID,
       PCIESS_AXI_1_S_AWADDR,
       PCIESS_AXI_1_S_AWBURST,
       PCIESS_AXI_1_S_AWID,
       PCIESS_AXI_1_S_AWLEN,
       PCIESS_AXI_1_S_AWSIZE,
       PCIESS_AXI_1_S_AWVALID,
       PCIESS_AXI_1_S_BREADY,
       PCIESS_AXI_1_S_RREADY,
       PCIESS_AXI_1_S_WLAST,
       PCIESS_AXI_1_S_WSTRB,
       PCIESS_AXI_1_S_WVALID,
       PCIE_1_TX_BIT_CLK,
       PCIE_1_TX_PLL_REF_CLK,
       PCIE_1_TX_PLL_LOCK,
       PCIESS_AXI_1_S_RDATA,
       PCIESS_AXI_1_S_WDATA,
       PCIESS_LANE2_CDR_REF_CLK_0,
       PCIESS_AXI_1_M_WDATA,
       PCIESS_AXI_1_M_RDATA
    );
output [31:0] APB_S_PRDATA;
output APB_S_PREADY;
output APB_S_PSLVERR;
input  [27:2] APB_S_PADDR;
input  APB_S_PENABLE;
input  APB_S_PSEL;
input  [31:0] APB_S_PWDATA;
input  APB_S_PWRITE;
input  APB_S_PCLK;
input  APB_S_PRESET_N;
input  PCIESS_LANE_RXD2_P;
input  PCIESS_LANE_RXD2_N;
output PCIESS_LANE_TXD2_P;
output PCIESS_LANE_TXD2_N;
input  AXI_CLK;
input  AXI_CLK_STABLE;
output [4:0] PCIE_1_LTSSM;
output PCIE_1_INTERRUPT_OUT;
input  [7:0] PCIE_1_INTERRUPT;
input  PCIE_1_TL_CLK_125MHz;
output PCIE_1_M_WDERR;
output PCIE_1_S_RDERR;
input  PCIE_1_M_RDERR;
input  PCIE_1_S_WDERR;
output PCIE_1_L2_EXIT;
output PCIE_1_HOT_RST_EXIT;
output PCIE_1_DLUP_EXIT;
input  PCIE_1_PERST_N;
output [3:0] PCIESS_AXI_1_M_ARID;
output [3:0] PCIESS_AXI_1_M_AWID;
output [31:0] PCIESS_AXI_1_M_ARADDR;
output [1:0] PCIESS_AXI_1_M_ARBURST;
output [7:0] PCIESS_AXI_1_M_ARLEN;
output [1:0] PCIESS_AXI_1_M_ARSIZE;
output PCIESS_AXI_1_M_ARVALID;
output [31:0] PCIESS_AXI_1_M_AWADDR;
output [1:0] PCIESS_AXI_1_M_AWBURST;
output [7:0] PCIESS_AXI_1_M_AWLEN;
output [1:0] PCIESS_AXI_1_M_AWSIZE;
output PCIESS_AXI_1_M_AWVALID;
output PCIESS_AXI_1_M_BREADY;
output PCIESS_AXI_1_M_RREADY;
output PCIESS_AXI_1_M_WLAST;
output [7:0] PCIESS_AXI_1_M_WSTRB;
output PCIESS_AXI_1_M_WVALID;
output PCIESS_AXI_1_S_ARREADY;
output PCIESS_AXI_1_S_AWREADY;
output [3:0] PCIESS_AXI_1_S_BID;
output [1:0] PCIESS_AXI_1_S_BRESP;
output PCIESS_AXI_1_S_BVALID;
output [3:0] PCIESS_AXI_1_S_RID;
output PCIESS_AXI_1_S_RLAST;
output [1:0] PCIESS_AXI_1_S_RRESP;
output PCIESS_AXI_1_S_RVALID;
output PCIESS_AXI_1_S_WREADY;
input  PCIESS_AXI_1_M_ARREADY;
input  PCIESS_AXI_1_M_AWREADY;
input  [3:0] PCIESS_AXI_1_M_BID;
input  [1:0] PCIESS_AXI_1_M_BRESP;
input  PCIESS_AXI_1_M_BVALID;
input  [3:0] PCIESS_AXI_1_M_RID;
input  PCIESS_AXI_1_M_RLAST;
input  [1:0] PCIESS_AXI_1_M_RRESP;
input  PCIESS_AXI_1_M_RVALID;
input  PCIESS_AXI_1_M_WREADY;
input  [31:0] PCIESS_AXI_1_S_ARADDR;
input  [1:0] PCIESS_AXI_1_S_ARBURST;
input  [3:0] PCIESS_AXI_1_S_ARID;
input  [7:0] PCIESS_AXI_1_S_ARLEN;
input  [1:0] PCIESS_AXI_1_S_ARSIZE;
input  PCIESS_AXI_1_S_ARVALID;
input  [31:0] PCIESS_AXI_1_S_AWADDR;
input  [1:0] PCIESS_AXI_1_S_AWBURST;
input  [3:0] PCIESS_AXI_1_S_AWID;
input  [7:0] PCIESS_AXI_1_S_AWLEN;
input  [1:0] PCIESS_AXI_1_S_AWSIZE;
input  PCIESS_AXI_1_S_AWVALID;
input  PCIESS_AXI_1_S_BREADY;
input  PCIESS_AXI_1_S_RREADY;
input  PCIESS_AXI_1_S_WLAST;
input  [7:0] PCIESS_AXI_1_S_WSTRB;
input  PCIESS_AXI_1_S_WVALID;
input  PCIE_1_TX_BIT_CLK;
input  PCIE_1_TX_PLL_REF_CLK;
input  PCIE_1_TX_PLL_LOCK;
output [63:0] PCIESS_AXI_1_S_RDATA;
input  [63:0] PCIESS_AXI_1_S_WDATA;
input  PCIESS_LANE2_CDR_REF_CLK_0;
output [63:0] PCIESS_AXI_1_M_WDATA;
input  [63:0] PCIESS_AXI_1_M_RDATA;

    wire 
        pcie_apblink_master_inst_lnk_m_rdata_pcie_apblink_inst_S_RDATA_net_0, 
        pcie_apblink_master_inst_lnk_m_rdata_pcie_apblink_inst_S_RDATA_net_1, 
        pcie_apblink_master_inst_lnk_m_rdata_pcie_apblink_inst_S_RDATA_net_2, 
        pcie_apblink_master_inst_lnk_m_rdata_pcie_apblink_inst_S_RDATA_net_3, 
        pcie_apblink_master_inst_lnk_m_rst_b_pcie_apblink_inst_S_ARST_N_net, 
        pcie_apblink_master_inst_lnk_m_enable_pcie_apblink_inst_S_EN_net, 
        pcie_apblink_master_inst_lnk_m_clock_pcie_apblink_inst_S_CLK_net, 
        pcie_apblink_master_inst_lnk_m_addr_pcie_apblink_inst_S_ADDR_net_0, 
        pcie_apblink_master_inst_lnk_m_addr_pcie_apblink_inst_S_ADDR_net_1, 
        pcie_apblink_master_inst_lnk_m_addr_pcie_apblink_inst_S_ADDR_net_2, 
        pcie_apblink_master_inst_lnk_m_wdata_pcie_apblink_inst_S_WDATA_net_0, 
        pcie_apblink_master_inst_lnk_m_wdata_pcie_apblink_inst_S_WDATA_net_1, 
        pcie_apblink_master_inst_lnk_m_wdata_pcie_apblink_inst_S_WDATA_net_2, 
        pcie_apblink_master_inst_lnk_m_wdata_pcie_apblink_inst_S_WDATA_net_3, 
        vcc_net, gnd_net, 
        pcie_apblink_inst_PCIE1_BRIDGE_CLK_PCIE_1_LINK_BRIDGE_CLK_net, 
        pcie_apblink_inst_PCIE1_BRIDGE_EN_PCIE_1_LINK_BRIDGE_EN_net, 
        pcie_apblink_inst_PCIE1_BRIDGE_ARST_N_PCIE_1_LINK_BRIDGE_ARST_N_net, 
        pcie_apblink_inst_PCIE1_BRIDGE_ADDR_PCIE_1_LINK_BRIDGE_ADDR_net_0, 
        pcie_apblink_inst_PCIE1_BRIDGE_ADDR_PCIE_1_LINK_BRIDGE_ADDR_net_1, 
        pcie_apblink_inst_PCIE1_BRIDGE_ADDR_PCIE_1_LINK_BRIDGE_ADDR_net_2, 
        pcie_apblink_inst_PCIE1_BRIDGE_RDATA_PCIE_1_LINK_BRIDGE_RDATA_net_0, 
        pcie_apblink_inst_PCIE1_BRIDGE_RDATA_PCIE_1_LINK_BRIDGE_RDATA_net_1, 
        pcie_apblink_inst_PCIE1_BRIDGE_RDATA_PCIE_1_LINK_BRIDGE_RDATA_net_2, 
        pcie_apblink_inst_PCIE1_BRIDGE_RDATA_PCIE_1_LINK_BRIDGE_RDATA_net_3, 
        pcie_apblink_inst_PCIE1_BRIDGE_WDATA_PCIE_1_LINK_BRIDGE_WDATA_net_0, 
        pcie_apblink_inst_PCIE1_BRIDGE_WDATA_PCIE_1_LINK_BRIDGE_WDATA_net_1, 
        pcie_apblink_inst_PCIE1_BRIDGE_WDATA_PCIE_1_LINK_BRIDGE_WDATA_net_2, 
        pcie_apblink_inst_PCIE1_BRIDGE_WDATA_PCIE_1_LINK_BRIDGE_WDATA_net_3, 
        PCIE_COMMON_AXI_CLK_OUT_net, 
        AXI_CLK_STABLE_FROM_PCIECOMMON_TO_PCIE_1_net, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_0, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_1, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_2, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_3, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_4, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_5, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_6, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_7, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_8, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_9, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_10, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_11, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_12, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_13, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_14, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_15, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_16, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_17, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_18, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_19, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_20, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_21, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_22, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_23, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_24, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_25, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_26, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_27, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_28, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_29, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_30, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_31, 
        PCIE_1_M_ARADDR_31_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_31_net, 
        PCIE_1_M_ARADDR_30_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_30_net, 
        PCIE_1_M_ARADDR_29_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_29_net, 
        PCIE_1_M_ARADDR_28_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_28_net, 
        PCIE_1_M_ARADDR_23_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_23_net, 
        PCIE_1_M_ARADDR_22_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_22_net, 
        PCIE_1_M_ARADDR_21_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_21_net, 
        PCIE_1_M_ARADDR_20_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_20_net, 
        PCIE_1_M_ARADDR_19_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_19_net, 
        PCIE_1_M_ARADDR_18_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_18_net, 
        PCIE_1_M_ARADDR_17_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_17_net, 
        PCIE_1_M_ARADDR_16_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_16_net, 
        PCIE_1_M_ARADDR_15_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_15_net, 
        PCIE_1_M_ARADDR_14_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_14_net, 
        PCIE_1_M_ARADDR_13_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_13_net, 
        PCIE_1_M_ARADDR_12_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_12_net, 
        PCIE_1_M_ARADDR_11_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_11_net, 
        PCIE_1_M_ARADDR_10_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_10_net, 
        PCIE_1_M_ARADDR_9_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_9_net, 
        PCIE_1_M_ARADDR_8_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_8_net, 
        PCIE_1_M_ARADDR_7_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_7_net, 
        PCIE_1_M_ARADDR_6_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_6_net, 
        PCIE_1_M_ARADDR_5_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_5_net, 
        PCIE_1_M_ARADDR_4_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_4_net, 
        PCIE_1_M_ARADDR_3_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_3_net, 
        PCIE_1_M_ARADDR_2_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_2_net, 
        PCIE_1_M_ARADDR_1_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_1_net, 
        PCIE_1_M_ARADDR_0_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_0_net, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_0, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_1, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_2, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_3, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_4, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_5, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_6, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_7, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_8, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_9, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_10, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_11, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_12, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_13, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_14, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_15, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_16, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_17, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_18, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_19, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_20, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_21, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_22, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_23, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_24, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_25, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_26, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_27, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_28, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_29, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_30, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_31, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_32, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_33, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_34, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_35, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_36, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_37, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_38, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_39, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_40, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_41, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_42, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_43, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_44, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_45, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_46, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_47, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_48, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_49, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_50, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_51, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_52, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_53, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_54, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_55, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_56, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_57, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_58, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_59, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_60, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_61, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_62, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_63, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_0, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_1, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_2, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_3, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_4, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_5, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_6, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_7, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_8, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_9, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_10, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_11, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_12, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_13, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_14, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_15, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_16, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_17, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_18, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_19, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_20, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_21, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_22, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_23, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_24, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_25, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_26, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_27, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_28, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_29, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_30, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_31, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_32, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_33, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_34, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_35, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_36, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_37, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_38, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_39, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_40, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_41, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_42, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_43, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_44, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_45, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_46, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_47, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_48, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_49, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_50, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_51, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_52, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_53, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_54, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_55, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_56, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_57, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_58, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_59, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_60, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_61, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_62, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_63, 
        PCIE_1_S_ARADDR_31_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_31_net, 
        PCIE_1_S_ARADDR_30_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_30_net, 
        PCIE_1_S_ARADDR_28_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_28_net, 
        PCIE_1_S_ARADDR_23_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_23_net, 
        PCIE_1_S_ARADDR_22_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_22_net, 
        PCIE_1_S_ARADDR_21_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_21_net, 
        PCIE_1_S_ARADDR_20_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_20_net, 
        PCIE_1_S_ARADDR_19_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_19_net, 
        PCIE_1_S_ARADDR_18_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_18_net, 
        PCIE_1_S_ARADDR_17_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_17_net, 
        PCIE_1_S_ARADDR_16_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_16_net, 
        PCIE_1_S_ARADDR_15_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_15_net, 
        PCIE_1_S_ARADDR_14_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_14_net, 
        PCIE_1_S_ARADDR_13_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_13_net, 
        PCIE_1_S_ARADDR_12_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_12_net, 
        PCIE_1_S_ARADDR_11_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_11_net, 
        PCIE_1_S_ARADDR_10_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_10_net, 
        PCIE_1_S_ARADDR_9_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_9_net, 
        PCIE_1_S_ARADDR_8_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_8_net, 
        PCIE_1_S_ARADDR_7_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_7_net, 
        PCIE_1_S_ARADDR_6_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_6_net, 
        PCIE_1_S_ARADDR_5_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_5_net, 
        PCIE_1_S_ARADDR_4_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_4_net, 
        PCIE_1_S_ARADDR_3_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_3_net, 
        PCIE_1_S_ARADDR_2_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_2_net, 
        PCIE_1_S_ARADDR_1_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_1_net, 
        PCIE_1_S_ARADDR_0_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_0_net, 
        PCIE_1_PHYSTATUS_2_PCIESS_LANE2_Pipe_AXI1_PHYSTATUS_0_net, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_0, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_1, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_2, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_3, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_4, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_5, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_6, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_7, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_8, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_9, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_10, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_11, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_12, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_13, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_14, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_15, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_16, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_17, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_18, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_19, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_20, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_21, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_22, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_23, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_24, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_25, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_26, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_27, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_28, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_29, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_30, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_31, 
        PCIE_1_RXDATAK_2_PCIESS_LANE2_Pipe_AXI1_RXDATAK_0_net_0, 
        PCIE_1_RXDATAK_2_PCIESS_LANE2_Pipe_AXI1_RXDATAK_0_net_1, 
        PCIE_1_RXDATAK_2_PCIESS_LANE2_Pipe_AXI1_RXDATAK_0_net_2, 
        PCIE_1_RXDATAK_2_PCIESS_LANE2_Pipe_AXI1_RXDATAK_0_net_3, 
        PCIE_1_RXELECIDLE_2_PCIESS_LANE2_Pipe_AXI1_RXELECIDLE_0_net, 
        PCIE_1_RXSTATUS_2_PCIESS_LANE2_Pipe_AXI1_RXSTATUS_0_net_0, 
        PCIE_1_RXSTATUS_2_PCIESS_LANE2_Pipe_AXI1_RXSTATUS_0_net_1, 
        PCIE_1_RXSTATUS_2_PCIESS_LANE2_Pipe_AXI1_RXSTATUS_0_net_2, 
        PCIE_1_RXVALID_2_PCIESS_LANE2_Pipe_AXI1_RXVALID_0_net, 
        PCIE_1_PCLK_OUT_2_PCIESS_LANE2_Pipe_AXI1_PCLK_OUT_0_net, 
        PCIE_1_RXPOLARITY_2_PCIESS_LANE2_Pipe_AXI1_RXPOLARITY_0_net, 
        PCIE_1_RXSTANDBYSTATUS_2_PCIESS_LANE2_Pipe_AXI1_RXSTANDBYSTATUS_0_net, 
        PCIE_1_TXCOMPLIANCE_2_PCIESS_LANE2_Pipe_AXI1_TXCOMPLIANCE_0_net, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_0, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_1, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_2, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_3, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_4, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_5, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_6, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_7, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_8, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_9, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_10, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_11, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_12, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_13, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_14, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_15, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_16, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_17, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_18, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_19, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_20, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_21, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_22, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_23, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_24, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_25, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_26, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_27, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_28, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_29, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_30, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_31, 
        PCIE_1_TXDATAK_2_PCIESS_LANE2_Pipe_AXI1_TXDATAK_0_net_0, 
        PCIE_1_TXDATAK_2_PCIESS_LANE2_Pipe_AXI1_TXDATAK_0_net_1, 
        PCIE_1_TXDATAK_2_PCIESS_LANE2_Pipe_AXI1_TXDATAK_0_net_2, 
        PCIE_1_TXDATAK_2_PCIESS_LANE2_Pipe_AXI1_TXDATAK_0_net_3, 
        PCIE_1_TXDATAVALID_2_PCIESS_LANE2_Pipe_AXI1_TXDATAVALID_0_net, 
        PCIE_1_TXDETECTRX_LOOPBACK_2_PCIESS_LANE2_Pipe_AXI1_TXDETECTRX_LOOPBACK_0_net, 
        PCIE_1_TXELECIDLE_2_PCIESS_LANE2_Pipe_AXI1_TXELECIDLE_0_net, 
        PCIE_1_PIPE_CLK_2_PCIESS_LANE2_Pipe_AXI1_PIPE_CLK_0_net, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_2_PCIESS_LANE2_Pipe_AXI1_PCS_DEBUG_net_0, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_2_PCIESS_LANE2_Pipe_AXI1_PCS_DEBUG_net_1, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_2_PCIESS_LANE2_Pipe_AXI1_PCS_DEBUG_net_2, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_2_PCIESS_LANE2_Pipe_AXI1_PCS_DEBUG_net_3, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_2_PCIESS_LANE2_Pipe_AXI1_PCS_DEBUG_net_4, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_2_PCIESS_LANE2_Pipe_AXI1_PCS_DEBUG_net_5, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_2_PCIESS_LANE2_Pipe_AXI1_PCS_DEBUG_net_6, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_2_PCIESS_LANE2_Pipe_AXI1_PCS_DEBUG_net_7, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_2_PCIESS_LANE2_Pipe_AXI1_PCS_DEBUG_net_8, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_2_PCIESS_LANE2_Pipe_AXI1_PCS_DEBUG_net_9, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_2_PCIESS_LANE2_Pipe_AXI1_PCS_DEBUG_net_10, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_2_PCIESS_LANE2_Pipe_AXI1_PCS_DEBUG_net_11, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_2_PCIESS_LANE2_Pipe_AXI1_PCS_DEBUG_net_12, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_2_PCIESS_LANE2_Pipe_AXI1_PCS_DEBUG_net_13, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_2_PCIESS_LANE2_Pipe_AXI1_PCS_DEBUG_net_14, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_2_PCIESS_LANE2_Pipe_AXI1_PCS_DEBUG_net_15, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_2_PCIESS_LANE2_Pipe_AXI1_PCS_DEBUG_net_16, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_2_PCIESS_LANE2_Pipe_AXI1_PCS_DEBUG_net_17, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_2_PCIESS_LANE2_Pipe_AXI1_PCS_DEBUG_net_18, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_2_PCIESS_LANE2_Pipe_AXI1_PCS_DEBUG_net_19, 
        PCIE_COMMON_INSTANCE_PMA_DEBUG_2_PCIESS_LANE2_Pipe_AXI1_PMA_DEBUG_net, 
        PCIE_1_M_AWADDR_31_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_31_net, 
        PCIE_1_M_AWADDR_30_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_30_net, 
        PCIE_1_M_AWADDR_29_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_29_net, 
        PCIE_1_M_AWADDR_28_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_28_net, 
        PCIE_1_M_AWADDR_23_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_23_net, 
        PCIE_1_M_AWADDR_22_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_22_net, 
        PCIE_1_M_AWADDR_21_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_21_net, 
        PCIE_1_M_AWADDR_20_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_20_net, 
        PCIE_1_M_AWADDR_19_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_19_net, 
        PCIE_1_M_AWADDR_18_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_18_net, 
        PCIE_1_M_AWADDR_17_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_17_net, 
        PCIE_1_M_AWADDR_16_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_16_net, 
        PCIE_1_M_AWADDR_15_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_15_net, 
        PCIE_1_M_AWADDR_14_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_14_net, 
        PCIE_1_M_AWADDR_13_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_13_net, 
        PCIE_1_M_AWADDR_12_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_12_net, 
        PCIE_1_M_AWADDR_11_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_11_net, 
        PCIE_1_M_AWADDR_10_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_10_net, 
        PCIE_1_M_AWADDR_9_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_9_net, 
        PCIE_1_M_AWADDR_8_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_8_net, 
        PCIE_1_M_AWADDR_7_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_7_net, 
        PCIE_1_M_AWADDR_6_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_6_net, 
        PCIE_1_M_AWADDR_5_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_5_net, 
        PCIE_1_M_AWADDR_4_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_4_net, 
        PCIE_1_M_AWADDR_3_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_3_net, 
        PCIE_1_M_AWADDR_2_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_2_net, 
        PCIE_1_M_AWADDR_1_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_1_net, 
        PCIE_1_M_AWADDR_0_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_0_net, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_0, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_1, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_2, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_3, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_4, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_5, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_6, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_7, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_8, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_9, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_10, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_11, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_12, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_13, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_14, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_15, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_16, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_17, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_18, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_19, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_20, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_21, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_22, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_23, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_24, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_25, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_26, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_27, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_28, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_29, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_30, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_31, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_32, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_33, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_34, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_35, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_36, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_37, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_38, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_39, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_40, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_41, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_42, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_43, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_44, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_45, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_46, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_47, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_48, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_49, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_50, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_51, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_52, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_53, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_54, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_55, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_56, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_57, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_58, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_59, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_60, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_61, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_62, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_63, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_0, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_1, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_2, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_3, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_4, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_5, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_6, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_7, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_8, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_9, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_10, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_11, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_12, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_13, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_14, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_15, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_16, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_17, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_18, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_19, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_20, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_21, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_22, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_23, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_24, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_25, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_26, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_27, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_28, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_29, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_30, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_31, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_32, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_33, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_34, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_35, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_36, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_37, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_38, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_39, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_40, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_41, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_42, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_43, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_44, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_45, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_46, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_47, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_48, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_49, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_50, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_51, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_52, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_53, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_54, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_55, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_56, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_57, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_58, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_59, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_60, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_61, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_62, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_63, 
        PCIE_1_S_AWADDR_31_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_31_net, 
        PCIE_1_S_AWADDR_30_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_30_net, 
        PCIE_1_S_AWADDR_28_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_28_net, 
        PCIE_1_S_AWADDR_23_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_23_net, 
        PCIE_1_S_AWADDR_22_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_22_net, 
        PCIE_1_S_AWADDR_21_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_21_net, 
        PCIE_1_S_AWADDR_20_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_20_net, 
        PCIE_1_S_AWADDR_19_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_19_net, 
        PCIE_1_S_AWADDR_18_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_18_net, 
        PCIE_1_S_AWADDR_17_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_17_net, 
        PCIE_1_S_AWADDR_16_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_16_net, 
        PCIE_1_S_AWADDR_15_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_15_net, 
        PCIE_1_S_AWADDR_14_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_14_net, 
        PCIE_1_S_AWADDR_13_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_13_net, 
        PCIE_1_S_AWADDR_12_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_12_net, 
        PCIE_1_S_AWADDR_11_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_11_net, 
        PCIE_1_S_AWADDR_10_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_10_net, 
        PCIE_1_S_AWADDR_9_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_9_net, 
        PCIE_1_S_AWADDR_8_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_8_net, 
        PCIE_1_S_AWADDR_7_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_7_net, 
        PCIE_1_S_AWADDR_6_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_6_net, 
        PCIE_1_S_AWADDR_5_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_5_net, 
        PCIE_1_S_AWADDR_4_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_4_net, 
        PCIE_1_S_AWADDR_3_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_3_net, 
        PCIE_1_S_AWADDR_2_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_2_net, 
        PCIE_1_S_AWADDR_1_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_1_net, 
        PCIE_1_S_AWADDR_0_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_0_net, 
        PCIE_1_PHYSTATUS_3_PCIESS_LANE3_Pipe_AXI0_PHYSTATUS_0_net, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_0, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_1, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_2, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_3, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_4, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_5, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_6, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_7, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_8, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_9, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_10, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_11, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_12, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_13, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_14, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_15, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_16, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_17, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_18, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_19, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_20, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_21, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_22, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_23, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_24, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_25, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_26, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_27, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_28, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_29, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_30, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_31, 
        PCIE_1_RXDATAK_3_PCIESS_LANE3_Pipe_AXI0_RXDATAK_0_net_0, 
        PCIE_1_RXDATAK_3_PCIESS_LANE3_Pipe_AXI0_RXDATAK_0_net_1, 
        PCIE_1_RXDATAK_3_PCIESS_LANE3_Pipe_AXI0_RXDATAK_0_net_2, 
        PCIE_1_RXDATAK_3_PCIESS_LANE3_Pipe_AXI0_RXDATAK_0_net_3, 
        PCIE_1_RXELECIDLE_3_PCIESS_LANE3_Pipe_AXI0_RXELECIDLE_0_net, 
        PCIE_1_RXSTATUS_3_PCIESS_LANE3_Pipe_AXI0_RXSTATUS_0_net_0, 
        PCIE_1_RXSTATUS_3_PCIESS_LANE3_Pipe_AXI0_RXSTATUS_0_net_1, 
        PCIE_1_RXSTATUS_3_PCIESS_LANE3_Pipe_AXI0_RXSTATUS_0_net_2, 
        PCIE_1_RXVALID_3_PCIESS_LANE3_Pipe_AXI0_RXVALID_0_net, 
        PCIE_1_PCLK_OUT_3_PCIESS_LANE3_Pipe_AXI0_PCLK_OUT_0_net, 
        PCIE_1_POWERDOWN_PCIESS_LANE2_Pipe_AXI1_POWERDOWN_net_0, 
        PCIE_1_POWERDOWN_PCIESS_LANE2_Pipe_AXI1_POWERDOWN_net_1, 
        PCIE_1_RATE_PCIESS_LANE2_Pipe_AXI1_RATE_net_0, 
        PCIE_1_RATE_PCIESS_LANE2_Pipe_AXI1_RATE_net_1, 
        PCIE_1_RESET_N_PCIESS_LANE2_Pipe_AXI1_RESET_N_net, 
        PCIE_1_RXPOLARITY_3_PCIESS_LANE3_Pipe_AXI0_RXPOLARITY_0_net, 
        PCIE_1_RXSTANDBYSTATUS_3_PCIESS_LANE3_Pipe_AXI0_RXSTANDBYSTATUS_0_net, 
        PCIE_1_TXCOMPLIANCE_3_PCIESS_LANE3_Pipe_AXI0_TXCOMPLIANCE_0_net, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_0, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_1, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_2, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_3, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_4, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_5, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_6, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_7, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_8, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_9, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_10, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_11, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_12, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_13, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_14, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_15, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_16, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_17, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_18, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_19, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_20, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_21, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_22, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_23, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_24, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_25, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_26, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_27, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_28, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_29, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_30, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_31, 
        PCIE_1_TXDATAK_3_PCIESS_LANE3_Pipe_AXI0_TXDATAK_0_net_0, 
        PCIE_1_TXDATAK_3_PCIESS_LANE3_Pipe_AXI0_TXDATAK_0_net_1, 
        PCIE_1_TXDATAK_3_PCIESS_LANE3_Pipe_AXI0_TXDATAK_0_net_2, 
        PCIE_1_TXDATAK_3_PCIESS_LANE3_Pipe_AXI0_TXDATAK_0_net_3, 
        PCIE_1_TXDATAVALID_3_PCIESS_LANE3_Pipe_AXI0_TXDATAVALID_0_net, 
        PCIE_1_TXDEEMPH_PCIESS_LANE2_Pipe_AXI1_TXDEEMPH_net, 
        PCIE_1_TXDETECTRX_LOOPBACK_3_PCIESS_LANE3_Pipe_AXI0_TXDETECTRX_LOOPBACK_0_net, 
        PCIE_1_TXELECIDLE_3_PCIESS_LANE3_Pipe_AXI0_TXELECIDLE_0_net, 
        PCIE_1_TXMARGIN_PCIESS_LANE2_Pipe_AXI1_TXMARGIN_net_0, 
        PCIE_1_TXMARGIN_PCIESS_LANE2_Pipe_AXI1_TXMARGIN_net_1, 
        PCIE_1_TXMARGIN_PCIESS_LANE2_Pipe_AXI1_TXMARGIN_net_2, 
        PCIE_1_TXSWING_PCIESS_LANE2_Pipe_AXI1_TXSWING_net, 
        PCIE_1_PIPE_CLK_3_PCIESS_LANE3_Pipe_AXI0_PIPE_CLK_0_net, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_3_PCIESS_LANE3_Pipe_AXI0_PCS_DEBUG_net_0, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_3_PCIESS_LANE3_Pipe_AXI0_PCS_DEBUG_net_1, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_3_PCIESS_LANE3_Pipe_AXI0_PCS_DEBUG_net_2, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_3_PCIESS_LANE3_Pipe_AXI0_PCS_DEBUG_net_3, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_3_PCIESS_LANE3_Pipe_AXI0_PCS_DEBUG_net_4, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_3_PCIESS_LANE3_Pipe_AXI0_PCS_DEBUG_net_5, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_3_PCIESS_LANE3_Pipe_AXI0_PCS_DEBUG_net_6, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_3_PCIESS_LANE3_Pipe_AXI0_PCS_DEBUG_net_7, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_3_PCIESS_LANE3_Pipe_AXI0_PCS_DEBUG_net_8, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_3_PCIESS_LANE3_Pipe_AXI0_PCS_DEBUG_net_9, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_3_PCIESS_LANE3_Pipe_AXI0_PCS_DEBUG_net_10, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_3_PCIESS_LANE3_Pipe_AXI0_PCS_DEBUG_net_11, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_3_PCIESS_LANE3_Pipe_AXI0_PCS_DEBUG_net_12, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_3_PCIESS_LANE3_Pipe_AXI0_PCS_DEBUG_net_13, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_3_PCIESS_LANE3_Pipe_AXI0_PCS_DEBUG_net_14, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_3_PCIESS_LANE3_Pipe_AXI0_PCS_DEBUG_net_15, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_3_PCIESS_LANE3_Pipe_AXI0_PCS_DEBUG_net_16, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_3_PCIESS_LANE3_Pipe_AXI0_PCS_DEBUG_net_17, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_3_PCIESS_LANE3_Pipe_AXI0_PCS_DEBUG_net_18, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_3_PCIESS_LANE3_Pipe_AXI0_PCS_DEBUG_net_19, 
        PCIE_COMMON_INSTANCE_PMA_DEBUG_3_PCIESS_LANE3_Pipe_AXI0_PMA_DEBUG_net;
    
    GND PCIESS_AXI_1_M_AWID_2_GndInst (.Y(PCIESS_AXI_1_M_AWID[2]));
    GND PCIESS_AXI_1_M_ARLEN_5_GndInst (.Y(PCIESS_AXI_1_M_ARLEN[5]));
    GND PCIESS_AXI_1_M_ARBURST_1_GndInst (.Y(PCIESS_AXI_1_M_ARBURST[1])
        );
    VCC vcc_inst (.Y(vcc_net));
    GND PCIESS_AXI_1_M_ARLEN_6_GndInst (.Y(PCIESS_AXI_1_M_ARLEN[6]));
    GND gnd_inst (.Y(gnd_net));
    GND PCIESS_AXI_1_M_AWLEN_7_GndInst (.Y(PCIESS_AXI_1_M_AWLEN[7]));
    PCIE_COMMON #( .MAIN_SOFT_RESET_NV_MAP(1'b0), .MAIN_SOFT_RESET_V_MAP(1'b0)
        , .MAIN_OVRLY_AXI0_IFC_MODE(2'b01), .MAIN_OVRLY_AXI1_IFC_MODE(2'b01)
        , .MAIN_INT_PIPE_CLK_CTRL_PCIE_0_PCLK_SEL(3'b110), .MAIN_INT_PIPE_CLK_CTRL_PCIE_1_PCLK_SEL(3'b010)
        , .MAIN_CLK_CTRL_AXI0_CLKENA(1'b0), .MAIN_CLK_CTRL_AXI1_CLKENA(1'b0)
        , .MAIN_DLL_STAT0_LOCK_INT_EN(1'b0), .MAIN_DLL_STAT0_UNLOCK_INT_EN(1'b0)
        , .MAIN_DLL_STAT0_LOCK_INT(1'b0), .MAIN_DLL_STAT0_UNLOCK_INT(1'b1)
        , .MAIN_TEST_DLL_RING_OSC_ENABLE(1'b0), .MAIN_TEST_DLL_REF_ENABLE(1'b0)
        , .MAIN_SPARE_SCRATCHPAD(8'b00000000), .MAIN_SPARE_SPARE_CTRL(24'b000000000000000000000000)
        , .MAIN_SOFT_RESET_PERIPH(1'b0), .MAIN_MAJOR_PCIE_USAGE_MODE(4'b1000)
        , .MAIN_INT_PIPE_CLK_CTRL_PCLK_INT_LN0_SEL(2'b10), .MAIN_INT_PIPE_CLK_CTRL_PCLK_INT_LN1_SEL(2'b10)
        , .MAIN_INT_PIPE_CLK_CTRL_PCLK_INT_LN2_SEL(1'b0), .MAIN_INT_PIPE_CLK_CTRL_PCLK_INT_LN3_SEL(1'b1)
        , .MAIN_EXT_PIPE_CLK_CTRL_PCLK_EXT_LN0_SEL(1'b0), .MAIN_EXT_PIPE_CLK_CTRL_PCLK_EXT_LN1_SEL(1'b0)
        , .MAIN_EXT_PIPE_CLK_CTRL_PCLK_EXT_LN2_SEL(1'b0), .MAIN_EXT_PIPE_CLK_CTRL_PCLK_EXT_LN3_SEL(1'b0)
        , .MAIN_QMUX_R0_PCIE_DBG_SEL(3'b111), .MAIN_DLL_CTRL0_PHASE_P(2'b11)
        , .MAIN_DLL_CTRL0_PHASE_S(2'b11), .MAIN_DLL_CTRL0_SEL_P(2'b00)
        , .MAIN_DLL_CTRL0_SEL_S(2'b00), .MAIN_DLL_CTRL0_REF_SEL(1'b0)
        , .MAIN_DLL_CTRL0_FB_SEL(1'b0), .MAIN_DLL_CTRL0_DIV_SEL(1'b0)
        , .MAIN_DLL_CTRL0_ALU_UPD(2'b00), .MAIN_DLL_CTRL0_LOCK_FRC(1'b0)
        , .MAIN_DLL_CTRL0_LOCK_FLT(2'b00), .MAIN_DLL_CTRL0_LOCK_HIGH(4'b1000)
        , .MAIN_DLL_CTRL0_LOCK_LOW(4'b1000), .MAIN_DLL_CTRL1_SET_ALU(8'b00000000)
        , .MAIN_DLL_CTRL1_ADJ_DEL4(7'b0000000), .MAIN_DLL_CTRL1_TEST_S(1'b0)
        , .MAIN_DLL_CTRL1_TEST_RING(1'b0), .MAIN_DLL_CTRL1_INIT_CODE(6'b000000)
        , .MAIN_DLL_CTRL1_RELOCK_FAST(1'b0), .MAIN_DLL_STAT0_RESET(1'b0)
        , .MAIN_DLL_STAT0_PHASE_MOVE_CLK(1'b0), .PMA_CMN_SOFT_RESET_PERIPH(1'b0)
        , .PCSCMN_SOFT_RESET_PERIPH(1'b0), .PCSCMN_GSSCLK_CTRL_MCLK_GSSCLK_0_SEL(5'b00000)
        , .PCSCMN_GSSCLK_CTRL_MCLK_GSSCLK_1_SEL(5'b00000), .PCSCMN_GSSCLK_CTRL_MCLK_GSSCLK_2_SEL(5'b00000)
        , .PCSCMN_QDBG_R0_PCS_DBG_MODE(3'b000), .PCSCMN_QDBG_R0_PCS_DBG_LANE_X(2'b00)
        , .PCSCMN_QDBG_R0_PCS_DBG_LANE_Y(2'b01) )  
        PCIE_COMMON_INSTANCE (.PHY_DEBUG({nc0, nc1, nc2, nc3}), 
        .PCS_DEBUG({nc4, nc5, nc6, nc7, nc8, nc9, nc10, nc11, nc12, 
        nc13, nc14, nc15, nc16, nc17, nc18, nc19, nc20, nc21, nc22, 
        nc23}), .PCIE_DEBUG({nc24, nc25, nc26, nc27, nc28, nc29, nc30, 
        nc31, nc32, nc33, nc34, nc35, nc36, nc37, nc38, nc39, nc40, 
        nc41, nc42, nc43, nc44, nc45, nc46, nc47, nc48, nc49, nc50, 
        nc51, nc52, nc53, nc54, nc55}), .AXI_CLK(AXI_CLK), 
        .AXI_CLK_STABLE(AXI_CLK_STABLE), .AXI_CLK_OUT(
        PCIE_COMMON_AXI_CLK_OUT_net), .PCS_DEBUG_0({gnd_net, gnd_net, 
        gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, 
        gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, 
        gnd_net, gnd_net, gnd_net, gnd_net}), .PMA_DEBUG_0(gnd_net), 
        .PCS_DEBUG_1({gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, 
        gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, 
        gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, 
        gnd_net}), .PMA_DEBUG_1(gnd_net), .PCS_DEBUG_2({
        PCIE_COMMON_INSTANCE_PCS_DEBUG_2_PCIESS_LANE2_Pipe_AXI1_PCS_DEBUG_net_19, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_2_PCIESS_LANE2_Pipe_AXI1_PCS_DEBUG_net_18, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_2_PCIESS_LANE2_Pipe_AXI1_PCS_DEBUG_net_17, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_2_PCIESS_LANE2_Pipe_AXI1_PCS_DEBUG_net_16, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_2_PCIESS_LANE2_Pipe_AXI1_PCS_DEBUG_net_15, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_2_PCIESS_LANE2_Pipe_AXI1_PCS_DEBUG_net_14, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_2_PCIESS_LANE2_Pipe_AXI1_PCS_DEBUG_net_13, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_2_PCIESS_LANE2_Pipe_AXI1_PCS_DEBUG_net_12, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_2_PCIESS_LANE2_Pipe_AXI1_PCS_DEBUG_net_11, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_2_PCIESS_LANE2_Pipe_AXI1_PCS_DEBUG_net_10, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_2_PCIESS_LANE2_Pipe_AXI1_PCS_DEBUG_net_9, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_2_PCIESS_LANE2_Pipe_AXI1_PCS_DEBUG_net_8, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_2_PCIESS_LANE2_Pipe_AXI1_PCS_DEBUG_net_7, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_2_PCIESS_LANE2_Pipe_AXI1_PCS_DEBUG_net_6, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_2_PCIESS_LANE2_Pipe_AXI1_PCS_DEBUG_net_5, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_2_PCIESS_LANE2_Pipe_AXI1_PCS_DEBUG_net_4, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_2_PCIESS_LANE2_Pipe_AXI1_PCS_DEBUG_net_3, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_2_PCIESS_LANE2_Pipe_AXI1_PCS_DEBUG_net_2, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_2_PCIESS_LANE2_Pipe_AXI1_PCS_DEBUG_net_1, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_2_PCIESS_LANE2_Pipe_AXI1_PCS_DEBUG_net_0})
        , .PMA_DEBUG_2(
        PCIE_COMMON_INSTANCE_PMA_DEBUG_2_PCIESS_LANE2_Pipe_AXI1_PMA_DEBUG_net)
        , .PCS_DEBUG_3({
        PCIE_COMMON_INSTANCE_PCS_DEBUG_3_PCIESS_LANE3_Pipe_AXI0_PCS_DEBUG_net_19, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_3_PCIESS_LANE3_Pipe_AXI0_PCS_DEBUG_net_18, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_3_PCIESS_LANE3_Pipe_AXI0_PCS_DEBUG_net_17, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_3_PCIESS_LANE3_Pipe_AXI0_PCS_DEBUG_net_16, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_3_PCIESS_LANE3_Pipe_AXI0_PCS_DEBUG_net_15, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_3_PCIESS_LANE3_Pipe_AXI0_PCS_DEBUG_net_14, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_3_PCIESS_LANE3_Pipe_AXI0_PCS_DEBUG_net_13, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_3_PCIESS_LANE3_Pipe_AXI0_PCS_DEBUG_net_12, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_3_PCIESS_LANE3_Pipe_AXI0_PCS_DEBUG_net_11, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_3_PCIESS_LANE3_Pipe_AXI0_PCS_DEBUG_net_10, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_3_PCIESS_LANE3_Pipe_AXI0_PCS_DEBUG_net_9, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_3_PCIESS_LANE3_Pipe_AXI0_PCS_DEBUG_net_8, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_3_PCIESS_LANE3_Pipe_AXI0_PCS_DEBUG_net_7, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_3_PCIESS_LANE3_Pipe_AXI0_PCS_DEBUG_net_6, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_3_PCIESS_LANE3_Pipe_AXI0_PCS_DEBUG_net_5, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_3_PCIESS_LANE3_Pipe_AXI0_PCS_DEBUG_net_4, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_3_PCIESS_LANE3_Pipe_AXI0_PCS_DEBUG_net_3, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_3_PCIESS_LANE3_Pipe_AXI0_PCS_DEBUG_net_2, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_3_PCIESS_LANE3_Pipe_AXI0_PCS_DEBUG_net_1, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_3_PCIESS_LANE3_Pipe_AXI0_PCS_DEBUG_net_0})
        , .PMA_DEBUG_3(
        PCIE_COMMON_INSTANCE_PMA_DEBUG_3_PCIESS_LANE3_Pipe_AXI0_PMA_DEBUG_net)
        , .PCIE_DEBUG_0({gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, 
        gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, 
        gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, 
        gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, 
        gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, gnd_net}), 
        .PCIE_DEBUG_1({
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_31, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_30, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_29, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_28, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_27, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_26, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_25, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_24, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_23, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_22, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_21, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_20, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_19, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_18, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_17, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_16, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_15, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_14, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_13, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_12, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_11, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_10, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_9, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_8, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_7, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_6, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_5, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_4, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_3, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_2, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_1, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_0}), 
        .DLL_OUT(), .AXI_CLK_STABLE_OUT(
        AXI_CLK_STABLE_FROM_PCIECOMMON_TO_PCIE_1_net));
    PCIE #( .MAIN_SOFT_RESET_PERIPH(1'b0), .MAIN_MAJOR_PCIE_USAGE_MODE(4'b1000)
        , .MAIN_INT_PIPE_CLK_CTRL_PCLK_INT_LN0_SEL(2'b10), .MAIN_INT_PIPE_CLK_CTRL_PCLK_INT_LN1_SEL(2'b10)
        , .MAIN_INT_PIPE_CLK_CTRL_PCLK_INT_LN2_SEL(1'b0), .MAIN_INT_PIPE_CLK_CTRL_PCLK_INT_LN3_SEL(1'b1)
        , .MAIN_EXT_PIPE_CLK_CTRL_PCLK_EXT_LN0_SEL(1'b0), .MAIN_EXT_PIPE_CLK_CTRL_PCLK_EXT_LN1_SEL(1'b0)
        , .MAIN_EXT_PIPE_CLK_CTRL_PCLK_EXT_LN2_SEL(1'b0), .MAIN_EXT_PIPE_CLK_CTRL_PCLK_EXT_LN3_SEL(1'b0)
        , .MAIN_QMUX_R0_PCIE_DBG_SEL(3'b111), .MAIN_DLL_CTRL0_PHASE_P(2'b11)
        , .MAIN_DLL_CTRL0_PHASE_S(2'b11), .MAIN_DLL_CTRL0_SEL_P(2'b00)
        , .MAIN_DLL_CTRL0_SEL_S(2'b00), .MAIN_DLL_CTRL0_REF_SEL(1'b0)
        , .MAIN_DLL_CTRL0_FB_SEL(1'b0), .MAIN_DLL_CTRL0_DIV_SEL(1'b0)
        , .MAIN_DLL_CTRL0_ALU_UPD(2'b00), .MAIN_DLL_CTRL0_LOCK_FRC(1'b0)
        , .MAIN_DLL_CTRL0_LOCK_FLT(2'b00), .MAIN_DLL_CTRL0_LOCK_HIGH(4'b1000)
        , .MAIN_DLL_CTRL0_LOCK_LOW(4'b1000), .MAIN_DLL_CTRL1_SET_ALU(8'b00000000)
        , .MAIN_DLL_CTRL1_ADJ_DEL4(7'b0000000), .MAIN_DLL_CTRL1_TEST_S(1'b0)
        , .MAIN_DLL_CTRL1_TEST_RING(1'b0), .MAIN_DLL_CTRL1_INIT_CODE(6'b000000)
        , .MAIN_DLL_CTRL1_RELOCK_FAST(1'b0), .MAIN_DLL_STAT0_RESET(1'b0)
        , .MAIN_DLL_STAT0_PHASE_MOVE_CLK(1'b0), .PMA_CMN_SOFT_RESET_PERIPH(1'b0)
        , .PCSCMN_SOFT_RESET_PERIPH(1'b0), .PCSCMN_GSSCLK_CTRL_MCLK_GSSCLK_0_SEL(5'b00000)
        , .PCSCMN_GSSCLK_CTRL_MCLK_GSSCLK_1_SEL(5'b00000), .PCSCMN_GSSCLK_CTRL_MCLK_GSSCLK_2_SEL(5'b00000)
        , .PCSCMN_QDBG_R0_PCS_DBG_MODE(3'b000), .PCSCMN_QDBG_R0_PCS_DBG_LANE_X(2'b00)
        , .PCSCMN_QDBG_R0_PCS_DBG_LANE_Y(2'b01), .PCSCMN_QRST_R0_QRST0_LANE(2'b00)
        , .PCSCMN_QRST_R0_QRST0_RST_SEL(4'b0000), .PCSCMN_QRST_R0_QRST1_LANE(2'b00)
        , .PCSCMN_QRST_R0_QRST1_RST_SEL(4'b0000), .MAIN_QMUX_R0_QRST0_SRC(3'b001)
        , .MAIN_QMUX_R0_QRST1_SRC(3'b011), .MAIN_QMUX_R0_QRST2_SRC(3'b000)
        , .MAIN_QMUX_R0_QRST3_SRC(3'b000), .PCIE_SITE("PCIE1"), .SIMULATION_MODE("BFM")
        , .REG_FILE(""), .MSC_UNIQUE(""), .SOFT_RESET_CTLR_CFG_BRGAXI_SOFTRST(1'b0)
        , .SOFT_RESET_CTLR_CFG_IGNORE_BRGAXI_SOFTRST_4_CTRL_RST(1'b1)
        , .SOFT_RESET_CTLR_CFG_IGNORE_MPERST(1'b0), .SOFT_RESET_CTLR_CFG_IGNORE_INBAND_RST_EVENT_4_CTRL_RST(1'b0)
        , .SOFT_RESET_CTLR_CFG_BRGMAP_SOFTRST(1'b0), .SOFT_RESET_CTLR_CFG_PCIE_CFGRESET_REL(1'b1)
        , .SEC_ERROR_INT_TX_RAM_SEC_ERR_INT(4'b0000), .SEC_ERROR_INT_RX_RAM_SEC_ERR_INT(4'b0000)
        , .SEC_ERROR_INT_PCIE2AXI_RAM_SEC_ERR_INT(4'b0000), .SEC_ERROR_INT_AXI2PCIE_RAM_SEC_ERR_INT(4'b0000)
        , .SEC_ERROR_INT_MASK_TX_RAM_SEC_ERR_INT_MASK(4'b0001), .SEC_ERROR_INT_MASK_RX_RAM_SEC_ERR_INT_MASK(4'b0001)
        , .SEC_ERROR_INT_MASK_PCIE2AXI_RAM_SEC_ERR_INT_MASK(4'b0001), .SEC_ERROR_INT_MASK_AXI2PCIE_RAM_SEC_ERR_INT_MASK(4'b0001)
        , .DED_ERROR_INT_TX_RAM_DED_ERR_INT(4'b0000), .DED_ERROR_INT_RX_RAM_DED_ERR_INT(4'b0000)
        , .DED_ERROR_INT_PCIE2AXI_RAM_DED_ERR_INT(4'b0000), .DED_ERROR_INT_AXI2PCIE_RAM_DED_ERR_INT(4'b0000)
        , .DED_ERROR_INT_MASK_TX_RAM_DED_ERR_INT_MASK(4'b0001), .DED_ERROR_INT_MASK_RX_RAM_DED_ERR_INT_MASK(4'b0001)
        , .DED_ERROR_INT_MASK_PCIE2AXI_RAM_DED_ERR_INT_MASK(4'b0001), .DED_ERROR_INT_MASK_AXI2PCIE_RAM_DED_ERR_INT_MASK(4'b0001)
        , .ECC_CONTROL_TX_RAM_INJ_ERR(4'b0000), .ECC_CONTROL_RX_RAM_INJ_ERR(4'b0000)
        , .ECC_CONTROL_PCIE2AXI_RAM_INJ_ERR(4'b0000), .ECC_CONTROL_AXI2PCIE_RAM_INJ_ERR(4'b0000)
        , .ECC_CONTROL_TX_RAM_ECC_BYPASS(1'b0), .ECC_CONTROL_RX_RAM_ECC_BYPASS(1'b0)
        , .ECC_CONTROL_PCIE2AXI_RAM_ECC_BYPASS(1'b0), .ECC_CONTROL_AXI2PCIE_RAM_ECC_BYPASS(1'b0)
        , .ECC_ERR_LOC_INJECT_ECC_ERR_ADDR(8'b00000000), .ECC_ERR_LOC_ENABLE_ECC_ERR_BIT_LOC(8'b00000000)
        , .ECC_ERR_LOC_ENABLE_ECC_ERR_BYTE_LOC(10'b0000000000), .RAM_MARGIN_1_RX_BUF_MARGIN(12'b000000000000)
        , .RAM_MARGIN_1_TX_BUF_MARGIN(12'b000000000000), .RAM_MARGIN_2_P2A_BUF_MARGIN(12'b000000000000)
        , .RAM_MARGIN_2_A2P_BUF_MARGIN(12'b000000000000), .RAM_POWER_CONTROL_RX_BUF_PWR_CTRL(3'b000)
        , .RAM_POWER_CONTROL_TX_BUF_PWR_CTRL(3'b000), .RAM_POWER_CONTROL_P2A_BUF_PWR_CTRL(3'b000)
        , .RAM_POWER_CONTROL_A2P_BUF_PWR_CTRL(3'b000), .DEBUG_SEL_FAB_DEBUG_SEL(8'b00000000)
        , .PL_WAKECLKREQ_PL_WAKE_OVERRIDE(1'b0), .PCIE_EVENT_INT_L2_EXIT_INT(1'b0)
        , .PCIE_EVENT_INT_HOTRST_EXIT_INT(1'b0), .PCIE_EVENT_INT_DLUP_EXIT_INT(1'b0)
        , .PCIE_EVENT_INT_L2_EXIT_INT_MASK(1'b0), .PCIE_EVENT_INT_HOTRST_EXIT_INT_MASK(1'b0)
        , .PCIE_EVENT_INT_DLUP_EXIT_INT_MASK(1'b0), .SPARE_SCRATCHPAD(8'b00000000)
        , .SPARE_SPARE_CTRL(24'b000000000000000000000000), .TEST_BUS_IN_31_0_TEST_BUS_IN_BIT0_SIM_MODE(1'b0)
        , .TEST_BUS_IN_31_0_TEST_BUS_IN_BIT1_DIS_LPWR_STATE_NEG(1'b0)
        , .TEST_BUS_IN_31_0_TEST_BUS_IN_BIT2_LBACK_MST(1'b0), .TEST_BUS_IN_31_0_TEST_BUS_IN_BIT3_EN_WARN_ASSERT(1'b0)
        , .TEST_BUS_IN_31_0_TEST_BUS_IN_BIT4_EN_INFO_ASSERT(1'b0), .TEST_BUS_IN_31_0_TEST_BUS_IN_BIT6_DIS_SCRAMBLING(1'b0)
        , .TEST_BUS_IN_31_0_TEST_BUS_IN_BIT7_CMPL_RCV_BIT(1'b0), .TEST_BUS_IN_31_0_TEST_BUS_IN_BIT8_TS2_DEEMPH_BIT_SEL(1'b0)
        , .TEST_BUS_IN_31_0_TEST_BUS_IN_BIT9_DIS_POLL_CMPL_ENTRY(1'b0)
        , .TEST_BUS_IN_31_0_TEST_BUS_IN_BIT10_FORCE_PLL_CMPL_ENTRY(1'b0)
        , .TEST_BUS_IN_31_0_TEST_BUS_IN_BIT14_DIS_PHY_STATUS_TO(1'b0)
        , .TEST_BUS_IN_31_0_TEST_BUS_IN_BIT18_NULLIFIED_WRTX(1'b0), .TEST_BUS_IN_31_0_TEST_BUS_IN_BIT19_EXT_SIM_MODE(1'b0)
        , .TEST_BUS_IN_31_0_TEST_BUS_IN_BIT20_CHECK_DCBALANCE(1'b0), .TEST_BUS_IN_31_0_TEST_BUS_IN_BIT21_DISABLE_SKP_PARITY(1'b0)
        , .TEST_BUS_IN_63_32_TEST_BUS_IN_BF_63_32(32'b00000000000000000000000000000000)
        , .BRIDGE_PCIE_BAR_01_DW0_BAR_SIZE_MASK(28'b1111111111111111000000000000)
        , .BRIDGE_PCIE_BAR_01_DW0_PREFETCH_OR_BAR_SIZE(1'b1), .BRIDGE_PCIE_BAR_01_DW0_ADDR_OR_BAR_SIZE(1'b1)
        , .BRIDGE_PCIE_BAR_01_DW0_BAR_TYPE(1'b0), .BRIDGE_PCIE_BAR_01_DW1_RESERVED_OR_BAR_SIZE_MASK(32'b11111111111111111111111111111111)
        , .BRIDGE_PCIE_BAR_23_DW0_BAR_SIZE_MASK(28'b1111111111110000000000000000)
        , .BRIDGE_PCIE_BAR_23_DW0_PREFETCH_OR_BAR_SIZE(1'b1), .BRIDGE_PCIE_BAR_23_DW0_ADDR_OR_BAR_SIZE(1'b1)
        , .BRIDGE_PCIE_BAR_23_DW0_BAR_TYPE(1'b0), .BRIDGE_PCIE_BAR_23_DW1_RESERVED_OR_BAR_SIZE_MASK(32'b11111111111111111111111111111111)
        , .BRIDGE_PCIE_BAR_45_DW0_BAR_SIZE_MASK(28'b0000000000000000000000000000)
        , .BRIDGE_PCIE_BAR_45_DW0_PREFETCH_OR_BAR_SIZE(1'b0), .BRIDGE_PCIE_BAR_45_DW0_ADDR_OR_BAR_SIZE(1'b0)
        , .BRIDGE_PCIE_BAR_45_DW0_BAR_TYPE(1'b0), .BRIDGE_PCIE_BAR_45_DW1_RESERVED_OR_BAR_SIZE_MASK(32'b00000000000000000000000000000000)
        , .BRIDGE_PCIE_BAR_WIN_PFETCH_MEMWIN_64BADDR(1'b0), .BRIDGE_PCIE_BAR_WIN_PFETCH_MEMWIN(1'b0)
        , .BRIDGE_PCIE_BAR_WIN_IOWIN_32BADDR(1'b0), .BRIDGE_PCIE_BAR_WIN_IOWIN(1'b0)
        , .BRIDGE_ATR0_PCIE_WIN0_SRCADDR_PARAM_SRC_ADDR_LDW(20'b00000000000000000000)
        , .BRIDGE_ATR0_PCIE_WIN0_SRCADDR_PARAM_ATR_SIZE(6'b001111), .BRIDGE_ATR0_PCIE_WIN0_SRCADDR_PARAM_ATR_IMPL(1'b1)
        , .BRIDGE_ATR0_PCIE_WIN0_SRC_ADDR_SRC_ADDR_UDW(32'b00000000000000000000000000000000)
        , .BRIDGE_ATR0_PCIE_WIN0_TRSL_ADDR_LSB_TRSL_ADDR_LDW(20'b00000011000000000000)
        , .BRIDGE_ATR0_PCIE_WIN0_TRSL_ADDR_UDW_TSLR_ADDR_UDW(32'b00000000000000000000000000000000)
        , .BRIDGE_ATR0_PCIE_WIN0_TRSL_PARAM_TRSF_PARAM(12'b000000000000)
        , .BRIDGE_ATR0_PCIE_WIN0_TRSL_PARAM_TRSL_ID(4'b0100), .BRIDGE_ATR1_PCIE_WIN0_SRCADDR_PARAM_SRC_ADDR_LDW(20'b00000000000000000000)
        , .BRIDGE_ATR1_PCIE_WIN0_SRCADDR_PARAM_ATR_SIZE(6'b001011), .BRIDGE_ATR1_PCIE_WIN0_SRCADDR_PARAM_ATR_IMPL(1'b0)
        , .BRIDGE_ATR1_PCIE_WIN0_SRC_ADDR_SRC_ADDR_UDW(32'b00000000000000000000000000000000)
        , .BRIDGE_ATR1_PCIE_WIN0_TRSL_ADDR_LSB_TRSL_ADDR_LDW(20'b00000000000000000000)
        , .BRIDGE_ATR1_PCIE_WIN0_TRSL_ADDR_UDW_TSLR_ADDR_UDW(32'b00000000000000000000000000000000)
        , .BRIDGE_ATR1_PCIE_WIN0_TRSL_PARAM_TRSF_PARAM(12'b000000000000)
        , .BRIDGE_ATR1_PCIE_WIN0_TRSL_PARAM_TRSL_ID(4'b0001), .BRIDGE_ATR2_PCIE_WIN0_SRCADDR_PARAM_SRC_ADDR_LDW(20'b00000000000000000000)
        , .BRIDGE_ATR2_PCIE_WIN0_SRCADDR_PARAM_ATR_SIZE(6'b010011), .BRIDGE_ATR2_PCIE_WIN0_SRCADDR_PARAM_ATR_IMPL(1'b1)
        , .BRIDGE_ATR2_PCIE_WIN0_SRC_ADDR_SRC_ADDR_UDW(32'b00000000000000000000000000000000)
        , .BRIDGE_ATR2_PCIE_WIN0_TRSL_ADDR_LSB_TRSL_ADDR_LDW(20'b00010000000000000000)
        , .BRIDGE_ATR2_PCIE_WIN0_TRSL_ADDR_UDW_TSLR_ADDR_UDW(32'b00000000000000000000000000000000)
        , .BRIDGE_ATR2_PCIE_WIN0_TRSL_PARAM_TRSF_PARAM(12'b000000000000)
        , .BRIDGE_ATR2_PCIE_WIN0_TRSL_PARAM_TRSL_ID(4'b0100), .BRIDGE_ATR3_PCIE_WIN0_SRCADDR_PARAM_SRC_ADDR_LDW(20'b00000000000000000000)
        , .BRIDGE_ATR3_PCIE_WIN0_SRCADDR_PARAM_ATR_SIZE(6'b001011), .BRIDGE_ATR3_PCIE_WIN0_SRCADDR_PARAM_ATR_IMPL(1'b0)
        , .BRIDGE_ATR3_PCIE_WIN0_SRC_ADDR_SRC_ADDR_UDW(32'b00000000000000000000000000000000)
        , .BRIDGE_ATR3_PCIE_WIN0_TRSL_ADDR_LSB_TRSL_ADDR_LDW(20'b00000000000000000000)
        , .BRIDGE_ATR3_PCIE_WIN0_TRSL_ADDR_UDW_TSLR_ADDR_UDW(32'b00000000000000000000000000000000)
        , .BRIDGE_ATR3_PCIE_WIN0_TRSL_PARAM_TRSF_PARAM(12'b000000000000)
        , .BRIDGE_ATR3_PCIE_WIN0_TRSL_PARAM_TRSL_ID(4'b0001), .BRIDGE_ATR4_PCIE_WIN0_SRCADDR_PARAM_SRC_ADDR_LDW(20'b00000000000000000000)
        , .BRIDGE_ATR4_PCIE_WIN0_SRCADDR_PARAM_ATR_SIZE(6'b001011), .BRIDGE_ATR4_PCIE_WIN0_SRCADDR_PARAM_ATR_IMPL(1'b0)
        , .BRIDGE_ATR4_PCIE_WIN0_SRC_ADDR_SRC_ADDR_UDW(32'b00000000000000000000000000000000)
        , .BRIDGE_ATR4_PCIE_WIN0_TRSL_ADDR_LSB_TRSL_ADDR_LDW(20'b00000000000000000000)
        , .BRIDGE_ATR4_PCIE_WIN0_TRSL_ADDR_UDW_TSLR_ADDR_UDW(32'b00000000000000000000000000000000)
        , .BRIDGE_ATR4_PCIE_WIN0_TRSL_PARAM_TRSF_PARAM(12'b000000000000)
        , .BRIDGE_ATR4_PCIE_WIN0_TRSL_PARAM_TRSL_ID(4'b0100), .BRIDGE_ATR5_PCIE_WIN0_SRCADDR_PARAM_SRC_ADDR_LDW(20'b00000000000000000000)
        , .BRIDGE_ATR5_PCIE_WIN0_SRCADDR_PARAM_ATR_SIZE(6'b001011), .BRIDGE_ATR5_PCIE_WIN0_SRCADDR_PARAM_ATR_IMPL(1'b0)
        , .BRIDGE_ATR5_PCIE_WIN0_SRC_ADDR_SRC_ADDR_UDW(32'b00000000000000000000000000000000)
        , .BRIDGE_ATR5_PCIE_WIN0_TRSL_ADDR_LSB_TRSL_ADDR_LDW(20'b00000000000000000000)
        , .BRIDGE_ATR5_PCIE_WIN0_TRSL_ADDR_UDW_TSLR_ADDR_UDW(32'b00000000000000000000000000000000)
        , .BRIDGE_ATR5_PCIE_WIN0_TRSL_PARAM_TRSF_PARAM(12'b000000000000)
        , .BRIDGE_ATR5_PCIE_WIN0_TRSL_PARAM_TRSL_ID(4'b0100), .BRIDGE_ATR0_PCIE_WIN1_SRCADDR_PARAM_SRC_ADDR_LDW(20'b00000000000000000000)
        , .BRIDGE_ATR0_PCIE_WIN1_SRCADDR_PARAM_ATR_SIZE(6'b001011), .BRIDGE_ATR0_PCIE_WIN1_SRCADDR_PARAM_ATR_IMPL(1'b0)
        , .BRIDGE_ATR0_PCIE_WIN1_SRC_ADDR_SRC_ADDR_UDW(32'b00000000000000000000000000000000)
        , .BRIDGE_ATR0_PCIE_WIN1_TRSL_ADDR_LSB_TRSL_ADDR_LDW(20'b00000000000000000000)
        , .BRIDGE_ATR0_PCIE_WIN1_TRSL_ADDR_UDW_TSLR_ADDR_UDW(32'b00000000000000000000000000000000)
        , .BRIDGE_ATR0_PCIE_WIN1_TRSL_PARAM_TRSF_PARAM(12'b000000000000)
        , .BRIDGE_ATR0_PCIE_WIN1_TRSL_PARAM_TRSL_ID(4'b1100), .BRIDGE_ATR1_PCIE_WIN1_SRCADDR_PARAM_SRC_ADDR_LDW(20'b00000000000000000000)
        , .BRIDGE_ATR1_PCIE_WIN1_SRCADDR_PARAM_ATR_SIZE(6'b001011), .BRIDGE_ATR1_PCIE_WIN1_SRCADDR_PARAM_ATR_IMPL(1'b0)
        , .BRIDGE_ATR1_PCIE_WIN1_SRC_ADDR_SRC_ADDR_UDW(32'b00000000000000000000000000000000)
        , .BRIDGE_ATR1_PCIE_WIN1_TRSL_ADDR_LSB_TRSL_ADDR_LDW(20'b00000000000000000000)
        , .BRIDGE_ATR1_PCIE_WIN1_TRSL_ADDR_UDW_TSLR_ADDR_UDW(32'b00000000000000000000000000000000)
        , .BRIDGE_ATR1_PCIE_WIN1_TRSL_PARAM_TRSF_PARAM(12'b000000000000)
        , .BRIDGE_ATR1_PCIE_WIN1_TRSL_PARAM_TRSL_ID(4'b0001), .BRIDGE_ATR2_PCIE_WIN1_SRCADDR_PARAM_SRC_ADDR_LDW(20'b00000000000000000000)
        , .BRIDGE_ATR2_PCIE_WIN1_SRCADDR_PARAM_ATR_SIZE(6'b001011), .BRIDGE_ATR2_PCIE_WIN1_SRCADDR_PARAM_ATR_IMPL(1'b0)
        , .BRIDGE_ATR2_PCIE_WIN1_SRC_ADDR_SRC_ADDR_UDW(32'b00000000000000000000000000000000)
        , .BRIDGE_ATR2_PCIE_WIN1_TRSL_ADDR_LSB_TRSL_ADDR_LDW(20'b00000000000000000000)
        , .BRIDGE_ATR2_PCIE_WIN1_TRSL_ADDR_UDW_TSLR_ADDR_UDW(32'b00000000000000000000000000000000)
        , .BRIDGE_ATR2_PCIE_WIN1_TRSL_PARAM_TRSF_PARAM(12'b000000000000)
        , .BRIDGE_ATR2_PCIE_WIN1_TRSL_PARAM_TRSL_ID(4'b0100), .BRIDGE_ATR3_PCIE_WIN1_SRCADDR_PARAM_SRC_ADDR_LDW(20'b00000000000000000000)
        , .BRIDGE_ATR3_PCIE_WIN1_SRCADDR_PARAM_ATR_SIZE(6'b001011), .BRIDGE_ATR3_PCIE_WIN1_SRCADDR_PARAM_ATR_IMPL(1'b0)
        , .BRIDGE_ATR3_PCIE_WIN1_SRC_ADDR_SRC_ADDR_UDW(32'b00000000000000000000000000000000)
        , .BRIDGE_ATR3_PCIE_WIN1_TRSL_ADDR_LSB_TRSL_ADDR_LDW(20'b00000000000000000000)
        , .BRIDGE_ATR3_PCIE_WIN1_TRSL_ADDR_UDW_TSLR_ADDR_UDW(32'b00000000000000000000000000000000)
        , .BRIDGE_ATR3_PCIE_WIN1_TRSL_PARAM_TRSF_PARAM(12'b000000000000)
        , .BRIDGE_ATR3_PCIE_WIN1_TRSL_PARAM_TRSL_ID(4'b0001), .BRIDGE_ATR4_PCIE_WIN1_SRCADDR_PARAM_SRC_ADDR_LDW(20'b00000000000000000000)
        , .BRIDGE_ATR4_PCIE_WIN1_SRCADDR_PARAM_ATR_SIZE(6'b001011), .BRIDGE_ATR4_PCIE_WIN1_SRCADDR_PARAM_ATR_IMPL(1'b0)
        , .BRIDGE_ATR4_PCIE_WIN1_SRC_ADDR_SRC_ADDR_UDW(32'b00000000000000000000000000000000)
        , .BRIDGE_ATR4_PCIE_WIN1_TRSL_ADDR_LSB_TRSL_ADDR_LDW(20'b00000000000000000000)
        , .BRIDGE_ATR4_PCIE_WIN1_TRSL_ADDR_UDW_TSLR_ADDR_UDW(32'b00000000000000000000000000000000)
        , .BRIDGE_ATR4_PCIE_WIN1_TRSL_PARAM_TRSF_PARAM(12'b000000000000)
        , .BRIDGE_ATR4_PCIE_WIN1_TRSL_PARAM_TRSL_ID(4'b0100), .BRIDGE_ATR5_PCIE_WIN1_SRCADDR_PARAM_SRC_ADDR_LDW(20'b00000000000000000000)
        , .BRIDGE_ATR5_PCIE_WIN1_SRCADDR_PARAM_ATR_SIZE(6'b001011), .BRIDGE_ATR5_PCIE_WIN1_SRCADDR_PARAM_ATR_IMPL(1'b0)
        , .BRIDGE_ATR5_PCIE_WIN1_SRC_ADDR_SRC_ADDR_UDW(32'b00000000000000000000000000000000)
        , .BRIDGE_ATR5_PCIE_WIN1_TRSL_ADDR_LSB_TRSL_ADDR_LDW(20'b00000000000000000000)
        , .BRIDGE_ATR5_PCIE_WIN1_TRSL_ADDR_UDW_TSLR_ADDR_UDW(32'b00000000000000000000000000000000)
        , .BRIDGE_ATR5_PCIE_WIN1_TRSL_PARAM_TRSF_PARAM(12'b000000000000)
        , .BRIDGE_ATR5_PCIE_WIN1_TRSL_PARAM_TRSL_ID(4'b0100), .BRIDGE_ATR0_AXI4_SLV0_SRCADDR_PARAM_SRC_ADDR_LDW(20'b00000000000000000000)
        , .BRIDGE_ATR0_AXI4_SLV0_SRCADDR_PARAM_ATR_SIZE(6'b001011), .BRIDGE_ATR0_AXI4_SLV0_SRCADDR_PARAM_ATR_IMPL(1'b0)
        , .BRIDGE_ATR0_AXI4_SLV0_SRC_ADDR_SRC_ADDR_UDW(32'b00000000000000000000000000000000)
        , .BRIDGE_ATR0_AXI4_SLV0_TRSL_ADDR_LSB_TRSL_ADDR_LDW(20'b00000000000000000000)
        , .BRIDGE_ATR0_AXI4_SLV0_TRSL_ADDR_UDW_TSLR_ADDR_UDW(32'b00000000000000000000000000000000)
        , .BRIDGE_ATR0_AXI4_SLV0_TRSL_PARAM_TRSF_PARAM(12'b000000000000)
        , .BRIDGE_ATR0_AXI4_SLV0_TRSL_PARAM_TRSL_ID(4'b0000), .BRIDGE_ATR1_AXI4_SLV0_SRCADDR_PARAM_SRC_ADDR_LDW(20'b00000000000000000000)
        , .BRIDGE_ATR1_AXI4_SLV0_SRCADDR_PARAM_ATR_SIZE(6'b001011), .BRIDGE_ATR1_AXI4_SLV0_SRCADDR_PARAM_ATR_IMPL(1'b0)
        , .BRIDGE_ATR1_AXI4_SLV0_SRC_ADDR_SRC_ADDR_UDW(32'b00000000000000000000000000000000)
        , .BRIDGE_ATR1_AXI4_SLV0_TRSL_ADDR_LSB_TRSL_ADDR_LDW(20'b00000000000000000000)
        , .BRIDGE_ATR1_AXI4_SLV0_TRSL_ADDR_UDW_TSLR_ADDR_UDW(32'b00000000000000000000000000000000)
        , .BRIDGE_ATR1_AXI4_SLV0_TRSL_PARAM_TRSF_PARAM(12'b000000000000)
        , .BRIDGE_ATR1_AXI4_SLV0_TRSL_PARAM_TRSL_ID(4'b0000), .BRIDGE_ATR2_AXI4_SLV0_SRCADDR_PARAM_SRC_ADDR_LDW(20'b00000000000000000000)
        , .BRIDGE_ATR2_AXI4_SLV0_SRCADDR_PARAM_ATR_SIZE(6'b001011), .BRIDGE_ATR2_AXI4_SLV0_SRCADDR_PARAM_ATR_IMPL(1'b0)
        , .BRIDGE_ATR2_AXI4_SLV0_SRC_ADDR_SRC_ADDR_UDW(32'b00000000000000000000000000000000)
        , .BRIDGE_ATR2_AXI4_SLV0_TRSL_ADDR_LSB_TRSL_ADDR_LDW(20'b00000000000000000000)
        , .BRIDGE_ATR2_AXI4_SLV0_TRSL_ADDR_UDW_TSLR_ADDR_UDW(32'b00000000000000000000000000000000)
        , .BRIDGE_ATR2_AXI4_SLV0_TRSL_PARAM_TRSF_PARAM(12'b000000000000)
        , .BRIDGE_ATR2_AXI4_SLV0_TRSL_PARAM_TRSL_ID(4'b0000), .BRIDGE_ATR3_AXI4_SLV0_SRCADDR_PARAM_SRC_ADDR_LDW(20'b00000000000000000000)
        , .BRIDGE_ATR3_AXI4_SLV0_SRCADDR_PARAM_ATR_SIZE(6'b001011), .BRIDGE_ATR3_AXI4_SLV0_SRCADDR_PARAM_ATR_IMPL(1'b0)
        , .BRIDGE_ATR3_AXI4_SLV0_SRC_ADDR_SRC_ADDR_UDW(32'b00000000000000000000000000000000)
        , .BRIDGE_ATR3_AXI4_SLV0_TRSL_ADDR_LSB_TRSL_ADDR_LDW(20'b00000000000000000000)
        , .BRIDGE_ATR3_AXI4_SLV0_TRSL_ADDR_UDW_TSLR_ADDR_UDW(32'b00000000000000000000000000000000)
        , .BRIDGE_ATR3_AXI4_SLV0_TRSL_PARAM_TRSF_PARAM(12'b000000000000)
        , .BRIDGE_ATR3_AXI4_SLV0_TRSL_PARAM_TRSL_ID(4'b0000), .BRIDGE_ATR4_AXI4_SLV0_SRCADDR_PARAM_SRC_ADDR_LDW(20'b00000000000000000000)
        , .BRIDGE_ATR4_AXI4_SLV0_SRCADDR_PARAM_ATR_SIZE(6'b001011), .BRIDGE_ATR4_AXI4_SLV0_SRCADDR_PARAM_ATR_IMPL(1'b0)
        , .BRIDGE_ATR4_AXI4_SLV0_SRC_ADDR_SRC_ADDR_UDW(32'b00000000000000000000000000000000)
        , .BRIDGE_ATR4_AXI4_SLV0_TRSL_ADDR_LSB_TRSL_ADDR_LDW(20'b00000000000000000000)
        , .BRIDGE_ATR4_AXI4_SLV0_TRSL_ADDR_UDW_TSLR_ADDR_UDW(32'b00000000000000000000000000000000)
        , .BRIDGE_ATR4_AXI4_SLV0_TRSL_PARAM_TRSF_PARAM(12'b000000000000)
        , .BRIDGE_ATR4_AXI4_SLV0_TRSL_PARAM_TRSL_ID(4'b0000), .BRIDGE_ATR5_AXI4_SLV0_SRCADDR_PARAM_SRC_ADDR_LDW(20'b00000000000000000000)
        , .BRIDGE_ATR5_AXI4_SLV0_SRCADDR_PARAM_ATR_SIZE(6'b001011), .BRIDGE_ATR5_AXI4_SLV0_SRCADDR_PARAM_ATR_IMPL(1'b0)
        , .BRIDGE_ATR5_AXI4_SLV0_SRC_ADDR_SRC_ADDR_UDW(32'b00000000000000000000000000000000)
        , .BRIDGE_ATR5_AXI4_SLV0_TRSL_ADDR_LSB_TRSL_ADDR_LDW(20'b00000000000000000000)
        , .BRIDGE_ATR5_AXI4_SLV0_TRSL_ADDR_UDW_TSLR_ADDR_UDW(32'b00000000000000000000000000000000)
        , .BRIDGE_ATR5_AXI4_SLV0_TRSL_PARAM_TRSF_PARAM(12'b000000000000)
        , .BRIDGE_ATR5_AXI4_SLV0_TRSL_PARAM_TRSL_ID(4'b0000), .BRIDGE_PCIE_VC_CRED_DW0_NP_DATA_CREDITS(4'b0000)
        , .BRIDGE_PCIE_VC_CRED_DW0_NP_HDR_CREDITS(8'b00010000), .BRIDGE_PCIE_VC_CRED_DW0_P_DATA_CREDITS(12'b000010111000)
        , .BRIDGE_PCIE_VC_CRED_DW0_P_HDR_CREDITS(8'b00011000), .BRIDGE_PCIE_VC_CRED_DW1_CPL_DATA_CREDITS(12'b000000000000)
        , .BRIDGE_PCIE_VC_CRED_DW1_CPL_HDR_CREDITS(8'b00000000), .BRIDGE_PCIE_VC_CRED_DW1_NP_DATA_CREDITS(4'b0001)
        , .BRIDGE_PCIE_PCI_IDS_DW0_DEVICE_ID(16'b0001010101010110), .BRIDGE_PCIE_PCI_IDS_DW0_VENDOR_ID(16'b0001000110101010)
        , .BRIDGE_PCIE_PCI_IDS_DW1_CLASS_CODE(24'b000000000000000000000000)
        , .BRIDGE_PCIE_PCI_IDS_DW1_REVISION_ID(8'b00000000), .BRIDGE_PCIE_PCI_IDS_DW2_SS_DEVICE_ID(16'b0000000000000000)
        , .BRIDGE_PCIE_PCI_IDS_DW2_SS_VENDOR_ID(16'b0000000000000000)
        , .BRIDGE_PCIE_PCI_LPM_PME_SUPPORT(5'b11111), .BRIDGE_PCIE_PCI_LPM_D2_SUPPORT(1'b1)
        , .BRIDGE_PCIE_PCI_LPM_D1_SUPPORT(1'b1), .BRIDGE_PCIE_PCI_LPM_AUX_CURRENT(3'b000)
        , .BRIDGE_PCIE_PCI_LPM_DSI(1'b0), .BRIDGE_PCIE_PCI_IRQ_DW0_MSIX_CAP(1'b1)
        , .BRIDGE_PCIE_PCI_IRQ_DW0_TABLE_SIZE(11'b00000000000), .BRIDGE_PCIE_PCI_IRQ_DW0_MSI_MASK_SUPPORT(1'b0)
        , .BRIDGE_PCIE_PCI_IRQ_DW0_NUM_MSI_MSGS(3'b010), .BRIDGE_PCIE_PCI_IRQ_DW0_INT_PIN(3'b100)
        , .BRIDGE_PCIE_PCI_IRQ_DW1_TABLE_OFFSET(29'b00000000000000000000000000000)
        , .BRIDGE_PCIE_PCI_IRQ_DW1_TABLE_BIR(3'b000), .BRIDGE_PCIE_PCI_IRQ_DW2_PBA_OFFSET(29'b00000000000000000000000000000)
        , .BRIDGE_PCIE_PCI_IRQ_DW2_PBA_BIR(3'b000), .BRIDGE_PCIE_PCI_IOV_DW0_ATS_PAGE_ALGN_REQ(1'b0)
        , .BRIDGE_PCIE_PCI_IOV_DW0_ATS_INVLD_QUEUE_DEPTH(5'b01010), .BRIDGE_PCIE_PCI_IOV_DW1_PRI_PAGE_REQ_CAP(32'b00000000000000000000000000000000)
        , .BRIDGE_PCIE_PEX_DEV_EP_L1_LATENCY(3'b000), .BRIDGE_PCIE_PEX_DEV_EP_L0_LATENCY(3'b000)
        , .BRIDGE_PCIE_PEX_DEV_MAXPAYLOAD(3'b001), .BRIDGE_PCIE_PEX_DEV2_LTR_SUPPORT(1'b1)
        , .BRIDGE_PCIE_PEX_DEV2_CPL_TIMEOUT_DISABLE(1'b1), .BRIDGE_PCIE_PEX_DEV2_CPL_TIMEOUT_RANGE(4'b1111)
        , .BRIDGE_PCIE_PEX_LINK_PORT_NUM(8'b00000001), .BRIDGE_PCIE_PEX_LINK_L1_EXIT_LATENCY(3'b000)
        , .BRIDGE_PCIE_PEX_LINK_L0S_EXIT_LATENCY(3'b001), .BRIDGE_PCIE_PEX_LINK_ASPM_L1(1'b1)
        , .BRIDGE_PCIE_PEX_LINK_ASPM_L0S(1'b1), .BRIDGE_PCIE_PEX_SPC_AER_IMPL(1'b1)
        , .BRIDGE_PCIE_PEX_SPC_DEV_NUM_RP(5'b00000), .BRIDGE_PCIE_PEX_SPC_RP_RCB(1'b0)
        , .BRIDGE_PCIE_PEX_SPC_LINK_SEL_DEEMPHASIS(1'b1), .BRIDGE_PCIE_PEX_SPC_SLOT_CLK_CFG(1'b0)
        , .BRIDGE_PCIE_PEX_SPC_SLOT_REG_IMPL(1'b1), .BRIDGE_PCIE_PEX_SPC2_ASPM_L1_DELAY(5'b00011)
        , .BRIDGE_PCIE_PEX_SPC2_ASPM_L0S_DELAY(5'b00011), .BRIDGE_PCIE_PEX_SPC2_PCIE_MSI_MSG_NUM(5'b00000)
        , .BRIDGE_PCIE_PEX_SPC2_AER_MSI_MSG_NUM(5'b00000), .BRIDGE_PCIE_PEX_SPC2_ECRC_CHK(1'b1)
        , .BRIDGE_PCIE_PEX_SPC2_ECRC_GEN(1'b1), .BRIDGE_PCIE_PEX_NFTS_NUM_FTS_8G(8'b00100000)
        , .BRIDGE_PCIE_PEX_NFTS_NUM_FTS_5G(8'b00100000), .BRIDGE_PCIE_PEX_NFTS_NUM_FTS_2P5G(8'b00100000)
        , .BRIDGE_PM_CONF_DW0_DATA_SCALE_7(2'b00), .BRIDGE_PM_CONF_DW0_DATA_SCALE_6(2'b00)
        , .BRIDGE_PM_CONF_DW0_DATA_SCALE_5(2'b00), .BRIDGE_PM_CONF_DW0_DATA_SCALE_4(2'b00)
        , .BRIDGE_PM_CONF_DW0_DATA_SCALE_3(2'b00), .BRIDGE_PM_CONF_DW0_DATA_SCALE_2(2'b00)
        , .BRIDGE_PM_CONF_DW0_DATA_SCALE_1(2'b00), .BRIDGE_PM_CONF_DW0_DATA_SCALE_0(2'b00)
        , .BRIDGE_PM_CONF_DW1_DATA_REGISTER_3(8'b00000000), .BRIDGE_PM_CONF_DW1_DATA_REGISTER_2(8'b00000000)
        , .BRIDGE_PM_CONF_DW1_DATA_REGISTER_1(8'b00000000), .BRIDGE_PM_CONF_DW1_DATA_REGISTER_0(8'b00000000)
        , .BRIDGE_PM_CONF_DW2_DATA_REGISTER_7(8'b00000000), .BRIDGE_PM_CONF_DW2_DATA_REGISTER_6(8'b00000000)
        , .BRIDGE_PM_CONF_DW2_DATA_REGISTER_5(8'b00000000), .BRIDGE_PM_CONF_DW2_DATA_REGISTER_4(8'b00000000)
        , .BRIDGE_PCIE_EQ_PRESET_DW0_UP_RCVR_PRST_LN1(3'b000), .BRIDGE_PCIE_EQ_PRESET_DW0_UP_XSMR_PRST_LN1(4'b0000)
        , .BRIDGE_PCIE_EQ_PRESET_DW0_DP_RCVR_PRST_LN1(3'b000), .BRIDGE_PCIE_EQ_PRESET_DW0_DP_XSMR_PRST_LN1(4'b0000)
        , .BRIDGE_PCIE_EQ_PRESET_DW0_UP_RCVR_PRST_LN0(3'b000), .BRIDGE_PCIE_EQ_PRESET_DW0_UP_XSMR_PRST_LN0(4'b0000)
        , .BRIDGE_PCIE_EQ_PRESET_DW0_DP_RCVR_PRST_LN0(3'b000), .BRIDGE_PCIE_EQ_PRESET_DW0_DP_XSMR_PRST_LN0(4'b0000)
        , .BRIDGE_PCIE_EQ_PRESET_DW1_UP_RCVR_PRST_LN3(3'b000), .BRIDGE_PCIE_EQ_PRESET_DW1_UP_XSMR_PRST_LN3(4'b0000)
        , .BRIDGE_PCIE_EQ_PRESET_DW1_DP_RCVR_PRST_LN3(3'b000), .BRIDGE_PCIE_EQ_PRESET_DW1_DP_XSMR_PRST_LN3(4'b0000)
        , .BRIDGE_PCIE_EQ_PRESET_DW1_UP_RCVR_PRST_LN2(3'b000), .BRIDGE_PCIE_EQ_PRESET_DW1_UP_XSMR_PRST_LN2(4'b0000)
        , .BRIDGE_PCIE_EQ_PRESET_DW1_DP_RCVR_PRST_LN2(3'b000), .BRIDGE_PCIE_EQ_PRESET_DW1_DP_XSMR_PRST_LN2(4'b0000)
        , .BRIDGE_PCIE_EQ_PRESET_DW2_UP_RCVR_PRST_LN5(3'b000), .BRIDGE_PCIE_EQ_PRESET_DW2_UP_XSMR_PRST_LN5(4'b0000)
        , .BRIDGE_PCIE_EQ_PRESET_DW2_DP_RCVR_PRST_LN5(3'b000), .BRIDGE_PCIE_EQ_PRESET_DW2_DP_XSMR_PRST_LN5(4'b0000)
        , .BRIDGE_PCIE_EQ_PRESET_DW2_UP_RCVR_PRST_LN4(3'b000), .BRIDGE_PCIE_EQ_PRESET_DW2_UP_XSMR_PRST_LN4(4'b0000)
        , .BRIDGE_PCIE_EQ_PRESET_DW2_DP_RCVR_PRST_LN4(3'b000), .BRIDGE_PCIE_EQ_PRESET_DW2_DP_XSMR_PRST_LN4(4'b0000)
        , .BRIDGE_PCIE_EQ_PRESET_DW3_UP_RCVR_PRST_LN7(3'b000), .BRIDGE_PCIE_EQ_PRESET_DW3_UP_XSMR_PRST_LN7(4'b0000)
        , .BRIDGE_PCIE_EQ_PRESET_DW3_DP_RCVR_PRST_LN7(3'b000), .BRIDGE_PCIE_EQ_PRESET_DW3_DP_XSMR_PRST_LN7(4'b0000)
        , .BRIDGE_PCIE_EQ_PRESET_DW3_UP_RCVR_PRST_LN6(3'b000), .BRIDGE_PCIE_EQ_PRESET_DW3_UP_XSMR_PRST_LN6(4'b0000)
        , .BRIDGE_PCIE_EQ_PRESET_DW3_DP_RCVR_PRST_LN6(3'b000), .BRIDGE_PCIE_EQ_PRESET_DW3_DP_XSMR_PRST_LN6(4'b0000)
        , .BRIDGE_PCIE_EQ_PRESET_DW4_UP_RCVR_PRST_LN9(3'b000), .BRIDGE_PCIE_EQ_PRESET_DW4_UP_XSMR_PRST_LN9(4'b0000)
        , .BRIDGE_PCIE_EQ_PRESET_DW4_DP_RCVR_PRST_LN9(3'b000), .BRIDGE_PCIE_EQ_PRESET_DW4_DP_XSMR_PRST_LN9(4'b0000)
        , .BRIDGE_PCIE_EQ_PRESET_DW4_UP_RCVR_PRST_LN8(3'b000), .BRIDGE_PCIE_EQ_PRESET_DW4_UP_XSMR_PRST_LN8(4'b0000)
        , .BRIDGE_PCIE_EQ_PRESET_DW4_DP_RCVR_PRST_LN8(3'b000), .BRIDGE_PCIE_EQ_PRESET_DW4_DP_XSMR_PRST_LN8(4'b0000)
        , .BRIDGE_PCIE_EQ_PRESET_DW5_UP_RCVR_PRST_LN11(3'b000), .BRIDGE_PCIE_EQ_PRESET_DW5_UP_XSMR_PRST_LN11(4'b0000)
        , .BRIDGE_PCIE_EQ_PRESET_DW5_DP_RCVR_PRST_LN11(3'b000), .BRIDGE_PCIE_EQ_PRESET_DW5_DP_XSMR_PRST_LN11(4'b0000)
        , .BRIDGE_PCIE_EQ_PRESET_DW5_UP_RCVR_PRST_LN10(3'b000), .BRIDGE_PCIE_EQ_PRESET_DW5_UP_XSMR_PRST_LN10(4'b0000)
        , .BRIDGE_PCIE_EQ_PRESET_DW5_DP_RCVR_PRST_LN10(3'b000), .BRIDGE_PCIE_EQ_PRESET_DW5_DP_XSMR_PRST_LN10(4'b0000)
        , .BRIDGE_PCIE_EQ_PRESET_DW6_UP_RCVR_PRST_LN13(3'b000), .BRIDGE_PCIE_EQ_PRESET_DW6_UP_XSMR_PRST_LN13(4'b0000)
        , .BRIDGE_PCIE_EQ_PRESET_DW6_DP_RCVR_PRST_LN13(3'b000), .BRIDGE_PCIE_EQ_PRESET_DW6_DP_XSMR_PRST_LN13(4'b0000)
        , .BRIDGE_PCIE_EQ_PRESET_DW6_UP_RCVR_PRST_LN12(3'b000), .BRIDGE_PCIE_EQ_PRESET_DW6_UP_XSMR_PRST_LN12(4'b0000)
        , .BRIDGE_PCIE_EQ_PRESET_DW6_DP_RCVR_PRST_LN12(3'b000), .BRIDGE_PCIE_EQ_PRESET_DW6_DP_XSMR_PRST_LN12(4'b0000)
        , .BRIDGE_PCIE_EQ_PRESET_DW7_UP_RCVR_PRST_LN15(3'b000), .BRIDGE_PCIE_EQ_PRESET_DW7_UP_XSMR_PRST_LN15(4'b0000)
        , .BRIDGE_PCIE_EQ_PRESET_DW7_DP_RCVR_PRST_LN15(3'b000), .BRIDGE_PCIE_EQ_PRESET_DW7_DP_XSMR_PRST_LN15(4'b0000)
        , .BRIDGE_PCIE_EQ_PRESET_DW7_UP_RCVR_PRST_LN14(3'b000), .BRIDGE_PCIE_EQ_PRESET_DW7_UP_XSMR_PRST_LN14(4'b0000)
        , .BRIDGE_PCIE_EQ_PRESET_DW7_DP_RCVR_PRST_LN14(3'b000), .BRIDGE_PCIE_EQ_PRESET_DW7_DP_XSMR_PRST_LN14(4'b0000)
        , .MAIN_OVRLY_AXI_IFC_MODE(2'b01), .MAIN_INT_PIPE_CLK_CTRL_PCLK_SEL(3'b010)
        , .MAIN_CLK_CTRL_AXI_CLKENA(1'b1), .DEV_CONTROL_ROOT_PORT_NEP(1'b0)
        , .DEV_CONTROL_LINK_WIDTH_X2_SUPPORT(1'b0), .DEV_CONTROL_LINK_WIDTH_X4_SUPPORT(1'b0)
        , .DEV_CONTROL_LINK_SPEED_5GBPS_SUPPORT(1'b1), .DEV_CONTROL_LANE_REVERSAL_SUPPORT(1'b1)
        , .DEV_CONTROL_USE_RXELECIDLE_TO_DETECT_ELECIDLE_ENTRY(1'b0), .DEV_CONTROL_ENABLE_NULLIFY_TLP_ON_TXBUF_ECC_ERR(1'b0)
        , .CLOCK_CONTROL_TL_CLOCK_FREQ(10'b0001111101), .PCICONF_PCI_IDS_OVERRIDE_PCICONF_OVERRIDE_EN(1'b0)
        , .PCICONF_PCI_IDS_31_0_PCI_VENDOR_ID(16'b0001000110101010), .PCICONF_PCI_IDS_31_0_PCI_DEVICE_ID(16'b0001010101010110)
        , .PCICONF_PCI_IDS_63_32_PCI_REVISION_ID(8'b00000000), .PCICONF_PCI_IDS_63_32_PCI_CLASS_CODE(24'b000000000000000000000000)
        , .PCICONF_PCI_IDS_95_64_PCI_SUBSYSTEM_VENDOR_ID(16'b0000000000000000)
        , .PCICONF_PCI_IDS_95_64_PCI_SUBSYSTEM_DEVICE_ID(16'b0000000000000000)
        , .PCIE_PEX_DEV_LINK_SPC2_PEX_DEV_LINK_SPC2_OVERRIDE_EN(1'b0)
        , .PCIE_PEX_DEV_LINK_SPC2_L0S_ENTRY_DELAY(5'b00000), .PCIE_PEX_DEV_LINK_SPC2_L0S_EXIT_DELAY(3'b000)
        , .PCIE_PEX_DEV_LINK_SPC2_L0S_ACC_LATENCY(3'b111), .PCIE_PEX_DEV_LINK_SPC2_L1_ENTRY_DELAY(5'b00000)
        , .PCIE_PEX_DEV_LINK_SPC2_L1_EXIT_DELAY(3'b000), .PCIE_PEX_DEV_LINK_SPC2_L1_ACC_LATENCY(3'b000)
        , .PCIE_PEX_SPC_PEX_SPC_OVERRIDE_EN(1'b0), .PCIE_PEX_SPC_PCIE_SLOT_CLK_CONF(1'b1)
        , .PCIE_PEX_SPC_PCIE_DE_EMPH_LVL(1'b0), .PCIE_AXI_MASTER_ATR_CFG0_PCIE_AXI_MASTER_ATR_OVERRIDE_EN(1'b0)
        , .PCIE_AXI_MASTER_ATR_CFG0_PCIE_AXI_MASTER_ATR_IMPL(1'b0), .PCIE_AXI_MASTER_ATR_CFG0_PCIE_AXI_MASTER_ATR_SIZE(6'b000000)
        , .PCIE_AXI_MASTER_ATR_CFG0_PCIE_AXI_MASTER_ATR_TRSL_ADDR_L(20'b00000000000000000000)
        , .PCIE_AXI_MASTER_ATR_CFG1_PCIE_AXI_MASTER_ATR_TRSL_ADDR_U(32'b00000000000000000000000000000000)
        , .PCIE_AXI_MASTER_ATR_CFG2_PCIE_AXI_MASTER_ATR_TRSL_ID(4'b0000)
        , .PCIE_AXI_MASTER_ATR_CFG2_PCIE_AXI_MASTER_ATR_TRSF_PARAM(12'b000000000000)
        , .AXI_SLAVE_PCIE_ATR_CFG0_AXI_SLAVE_PCIE_ATR_OVERRIDE_EN(1'b0)
        , .AXI_SLAVE_PCIE_ATR_CFG0_AXI_SLAVE_PCIE_ATR_IMPL(1'b0), .AXI_SLAVE_PCIE_ATR_CFG0_AXI_SLAVE_PCIE_ATR_SIZE(6'b000000)
        , .AXI_SLAVE_PCIE_ATR_CFG0_AXI_SLAVE_PCIE_ATR_TRSL_ADDR_L(20'b00000000000000000000)
        , .AXI_SLAVE_PCIE_ATR_CFG1_AXI_SLAVE_PCIE_ATR_TRSL_ADDR_U(32'b00000000000000000000000000000000)
        , .AXI_SLAVE_PCIE_ATR_CFG2_AXI_SLAVE_PCIE_ATR_TRSL_ID(4'b0000)
        , .AXI_SLAVE_PCIE_ATR_CFG2_AXI_SLAVE_PCIE_ATR_TRSF_PARAM(12'b000000000000)
        , .PCIE_BAR_01_PEX_BAR01_OVERRIDE_EN(1'b0), .PCIE_BAR_01_PEX_BAR0_CTRL(4'b0000)
        , .PCIE_BAR_01_PEX_BAR0_SIZE(5'b00000), .PCIE_BAR_01_PEX_BAR1_CTRL(4'b0000)
        , .PCIE_BAR_01_PEX_BAR1_SIZE(5'b00000), .PCIE_BAR_23_PEX_BAR23_OVERRIDE_EN(1'b0)
        , .PCIE_BAR_23_PEX_BAR2_CTRL(4'b0000), .PCIE_BAR_23_PEX_BAR2_SIZE(5'b00000)
        , .PCIE_BAR_23_PEX_BAR3_CTRL(4'b0000), .PCIE_BAR_23_PEX_BAR3_SIZE(5'b00000)
        , .PCIE_BAR_45_PEX_BAR45_OVERRIDE_EN(1'b0), .PCIE_BAR_45_PEX_BAR4_CTRL(4'b0000)
        , .PCIE_BAR_45_PEX_BAR4_SIZE(5'b00000), .PCIE_BAR_45_PEX_BAR5_CTRL(4'b0000)
        , .PCIE_BAR_45_PEX_BAR5_SIZE(5'b00000), .PCIE_BAR_WIN_PEX_BAR_WIN_OVERRIDE_EN(1'b0)
        , .PCIE_BAR_WIN_PEX_BAR_WIN_CTRL(4'b0000) )  PCIE_1 (
        .M_ARADDR_24(PCIESS_AXI_1_M_ARADDR[24]), .M_ARADDR_25(
        PCIESS_AXI_1_M_ARADDR[25]), .M_ARADDR_26(
        PCIESS_AXI_1_M_ARADDR[26]), .M_ARADDR_27(
        PCIESS_AXI_1_M_ARADDR[27]), .M_ARBURST({nc56, 
        PCIESS_AXI_1_M_ARBURST[0]}), .M_ARID({PCIESS_AXI_1_M_ARID[3], 
        PCIESS_AXI_1_M_ARID[2], PCIESS_AXI_1_M_ARID[1], 
        PCIESS_AXI_1_M_ARID[0]}), .M_ARLEN({nc57, nc58, nc59, 
        PCIESS_AXI_1_M_ARLEN[4], PCIESS_AXI_1_M_ARLEN[3], 
        PCIESS_AXI_1_M_ARLEN[2], PCIESS_AXI_1_M_ARLEN[1], 
        PCIESS_AXI_1_M_ARLEN[0]}), .M_ARSIZE({PCIESS_AXI_1_M_ARSIZE[1], 
        PCIESS_AXI_1_M_ARSIZE[0]}), .M_ARVALID(PCIESS_AXI_1_M_ARVALID), 
        .M_AWADDR_24(PCIESS_AXI_1_M_AWADDR[24]), .M_AWADDR_25(
        PCIESS_AXI_1_M_AWADDR[25]), .M_AWADDR_26(
        PCIESS_AXI_1_M_AWADDR[26]), .M_AWADDR_27(
        PCIESS_AXI_1_M_AWADDR[27]), .M_AWBURST({nc60, 
        PCIESS_AXI_1_M_AWBURST[0]}), .M_AWID({nc61, nc62, 
        PCIESS_AXI_1_M_AWID[1], PCIESS_AXI_1_M_AWID[0]}), .M_AWLEN({
        nc63, nc64, nc65, PCIESS_AXI_1_M_AWLEN[4], 
        PCIESS_AXI_1_M_AWLEN[3], PCIESS_AXI_1_M_AWLEN[2], 
        PCIESS_AXI_1_M_AWLEN[1], PCIESS_AXI_1_M_AWLEN[0]}), .M_AWSIZE({
        PCIESS_AXI_1_M_AWSIZE[1], PCIESS_AXI_1_M_AWSIZE[0]}), 
        .M_AWVALID(PCIESS_AXI_1_M_AWVALID), .M_BREADY(
        PCIESS_AXI_1_M_BREADY), .M_RREADY(PCIESS_AXI_1_M_RREADY), 
        .M_WDERR(PCIE_1_M_WDERR), .M_WLAST(PCIESS_AXI_1_M_WLAST), 
        .M_WSTRB({PCIESS_AXI_1_M_WSTRB[7], PCIESS_AXI_1_M_WSTRB[6], 
        PCIESS_AXI_1_M_WSTRB[5], PCIESS_AXI_1_M_WSTRB[4], 
        PCIESS_AXI_1_M_WSTRB[3], PCIESS_AXI_1_M_WSTRB[2], 
        PCIESS_AXI_1_M_WSTRB[1], PCIESS_AXI_1_M_WSTRB[0]}), .M_WVALID(
        PCIESS_AXI_1_M_WVALID), .S_ARREADY(PCIESS_AXI_1_S_ARREADY), 
        .S_AWREADY(PCIESS_AXI_1_S_AWREADY), .S_BID({
        PCIESS_AXI_1_S_BID[3], PCIESS_AXI_1_S_BID[2], 
        PCIESS_AXI_1_S_BID[1], PCIESS_AXI_1_S_BID[0]}), .S_BRESP({
        PCIESS_AXI_1_S_BRESP[1], PCIESS_AXI_1_S_BRESP[0]}), .S_BVALID(
        PCIESS_AXI_1_S_BVALID), .S_RDERR(PCIE_1_S_RDERR), .S_RID({
        PCIESS_AXI_1_S_RID[3], PCIESS_AXI_1_S_RID[2], 
        PCIESS_AXI_1_S_RID[1], PCIESS_AXI_1_S_RID[0]}), .S_RLAST(
        PCIESS_AXI_1_S_RLAST), .S_RRESP({PCIESS_AXI_1_S_RRESP[1], 
        PCIESS_AXI_1_S_RRESP[0]}), .S_RVALID(PCIESS_AXI_1_S_RVALID), 
        .S_WREADY(PCIESS_AXI_1_S_WREADY), .L2_EXIT(PCIE_1_L2_EXIT), 
        .HOT_RST_EXIT(PCIE_1_HOT_RST_EXIT), .DLUP_EXIT(
        PCIE_1_DLUP_EXIT), .INTERRUPT_OUT(PCIE_1_INTERRUPT_OUT), 
        .LTSSM({PCIE_1_LTSSM[4], PCIE_1_LTSSM[3], PCIE_1_LTSSM[2], 
        PCIE_1_LTSSM[1], PCIE_1_LTSSM[0]}), .WAKEREQ_OEN(), .M_ARREADY(
        PCIESS_AXI_1_M_ARREADY), .M_AWREADY(PCIESS_AXI_1_M_AWREADY), 
        .M_BID({PCIESS_AXI_1_M_BID[3], PCIESS_AXI_1_M_BID[2], 
        PCIESS_AXI_1_M_BID[1], PCIESS_AXI_1_M_BID[0]}), .M_BRESP({
        PCIESS_AXI_1_M_BRESP[1], PCIESS_AXI_1_M_BRESP[0]}), .M_BVALID(
        PCIESS_AXI_1_M_BVALID), .M_RDERR(PCIE_1_M_RDERR), .M_RID({
        PCIESS_AXI_1_M_RID[3], PCIESS_AXI_1_M_RID[2], 
        PCIESS_AXI_1_M_RID[1], PCIESS_AXI_1_M_RID[0]}), .M_RLAST(
        PCIESS_AXI_1_M_RLAST), .M_RRESP({PCIESS_AXI_1_M_RRESP[1], 
        PCIESS_AXI_1_M_RRESP[0]}), .M_RVALID(PCIESS_AXI_1_M_RVALID), 
        .M_WREADY(PCIESS_AXI_1_M_WREADY), .S_ARADDR_24(
        PCIESS_AXI_1_S_ARADDR[24]), .S_ARADDR_25(
        PCIESS_AXI_1_S_ARADDR[25]), .S_ARADDR_26(
        PCIESS_AXI_1_S_ARADDR[26]), .S_ARADDR_27(
        PCIESS_AXI_1_S_ARADDR[27]), .S_ARADDR_29(
        PCIESS_AXI_1_S_ARADDR[29]), .S_ARBURST({
        PCIESS_AXI_1_S_ARBURST[1], PCIESS_AXI_1_S_ARBURST[0]}), 
        .S_ARID({PCIESS_AXI_1_S_ARID[3], PCIESS_AXI_1_S_ARID[2], 
        PCIESS_AXI_1_S_ARID[1], PCIESS_AXI_1_S_ARID[0]}), .S_ARLEN({
        PCIESS_AXI_1_S_ARLEN[7], PCIESS_AXI_1_S_ARLEN[6], 
        PCIESS_AXI_1_S_ARLEN[5], PCIESS_AXI_1_S_ARLEN[4], 
        PCIESS_AXI_1_S_ARLEN[3], PCIESS_AXI_1_S_ARLEN[2], 
        PCIESS_AXI_1_S_ARLEN[1], PCIESS_AXI_1_S_ARLEN[0]}), .S_ARSIZE({
        PCIESS_AXI_1_S_ARSIZE[1], PCIESS_AXI_1_S_ARSIZE[0]}), 
        .S_ARVALID(PCIESS_AXI_1_S_ARVALID), .S_AWADDR_24(
        PCIESS_AXI_1_S_AWADDR[24]), .S_AWADDR_25(
        PCIESS_AXI_1_S_AWADDR[25]), .S_AWADDR_26(
        PCIESS_AXI_1_S_AWADDR[26]), .S_AWADDR_27(
        PCIESS_AXI_1_S_AWADDR[27]), .S_AWADDR_29(
        PCIESS_AXI_1_S_AWADDR[29]), .S_AWBURST({
        PCIESS_AXI_1_S_AWBURST[1], PCIESS_AXI_1_S_AWBURST[0]}), 
        .S_AWID({PCIESS_AXI_1_S_AWID[3], PCIESS_AXI_1_S_AWID[2], 
        PCIESS_AXI_1_S_AWID[1], PCIESS_AXI_1_S_AWID[0]}), .S_AWLEN({
        gnd_net, gnd_net, gnd_net, PCIESS_AXI_1_S_AWLEN[4], 
        PCIESS_AXI_1_S_AWLEN[3], PCIESS_AXI_1_S_AWLEN[2], 
        PCIESS_AXI_1_S_AWLEN[1], PCIESS_AXI_1_S_AWLEN[0]}), .S_AWSIZE({
        PCIESS_AXI_1_S_AWSIZE[1], PCIESS_AXI_1_S_AWSIZE[0]}), 
        .S_AWVALID(PCIESS_AXI_1_S_AWVALID), .S_BREADY(
        PCIESS_AXI_1_S_BREADY), .S_RREADY(PCIESS_AXI_1_S_RREADY), 
        .S_WDERR(PCIE_1_S_WDERR), .S_WLAST(PCIESS_AXI_1_S_WLAST), 
        .S_WSTRB({PCIESS_AXI_1_S_WSTRB[7], PCIESS_AXI_1_S_WSTRB[6], 
        PCIESS_AXI_1_S_WSTRB[5], PCIESS_AXI_1_S_WSTRB[4], 
        PCIESS_AXI_1_S_WSTRB[3], PCIESS_AXI_1_S_WSTRB[2], 
        PCIESS_AXI_1_S_WSTRB[1], PCIESS_AXI_1_S_WSTRB[0]}), .S_WVALID(
        PCIESS_AXI_1_S_WVALID), .INTERRUPT({PCIE_1_INTERRUPT[7], 
        PCIE_1_INTERRUPT[6], PCIE_1_INTERRUPT[5], PCIE_1_INTERRUPT[4], 
        PCIE_1_INTERRUPT[3], PCIE_1_INTERRUPT[2], PCIE_1_INTERRUPT[1], 
        PCIE_1_INTERRUPT[0]}), .MPERST_N(PCIE_1_PERST_N), .TL_CLK(
        PCIE_1_TL_CLK_125MHz), .WAKEREQ(vcc_net), .M_ARADDR_31(
        PCIE_1_M_ARADDR_31_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_31_net), 
        .M_ARADDR_30(
        PCIE_1_M_ARADDR_30_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_30_net), 
        .M_ARADDR_29(
        PCIE_1_M_ARADDR_29_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_29_net), 
        .M_ARADDR_28(
        PCIE_1_M_ARADDR_28_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_28_net), 
        .M_ARADDR_0(
        PCIE_1_M_ARADDR_0_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_0_net), 
        .M_ARADDR_1(
        PCIE_1_M_ARADDR_1_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_1_net), 
        .M_ARADDR_2(
        PCIE_1_M_ARADDR_2_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_2_net), 
        .M_ARADDR_3(
        PCIE_1_M_ARADDR_3_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_3_net), 
        .M_ARADDR_4(
        PCIE_1_M_ARADDR_4_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_4_net), 
        .M_ARADDR_5(
        PCIE_1_M_ARADDR_5_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_5_net), 
        .M_ARADDR_6(
        PCIE_1_M_ARADDR_6_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_6_net), 
        .M_ARADDR_7(
        PCIE_1_M_ARADDR_7_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_7_net), 
        .M_ARADDR_8(
        PCIE_1_M_ARADDR_8_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_8_net), 
        .M_ARADDR_9(
        PCIE_1_M_ARADDR_9_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_9_net), 
        .M_ARADDR_10(
        PCIE_1_M_ARADDR_10_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_10_net), 
        .M_ARADDR_11(
        PCIE_1_M_ARADDR_11_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_11_net), 
        .M_ARADDR_12(
        PCIE_1_M_ARADDR_12_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_12_net), 
        .M_ARADDR_13(
        PCIE_1_M_ARADDR_13_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_13_net), 
        .M_ARADDR_14(
        PCIE_1_M_ARADDR_14_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_14_net), 
        .M_ARADDR_15(
        PCIE_1_M_ARADDR_15_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_15_net), 
        .M_ARADDR_16(
        PCIE_1_M_ARADDR_16_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_16_net), 
        .M_ARADDR_17(
        PCIE_1_M_ARADDR_17_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_17_net), 
        .M_ARADDR_18(
        PCIE_1_M_ARADDR_18_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_18_net), 
        .M_ARADDR_19(
        PCIE_1_M_ARADDR_19_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_19_net), 
        .M_ARADDR_20(
        PCIE_1_M_ARADDR_20_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_20_net), 
        .M_ARADDR_21(
        PCIE_1_M_ARADDR_21_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_21_net), 
        .M_ARADDR_22(
        PCIE_1_M_ARADDR_22_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_22_net), 
        .M_ARADDR_23(
        PCIE_1_M_ARADDR_23_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_23_net), 
        .M_AWADDR_31(
        PCIE_1_M_AWADDR_31_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_31_net), 
        .M_AWADDR_30(
        PCIE_1_M_AWADDR_30_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_30_net), 
        .M_AWADDR_29(
        PCIE_1_M_AWADDR_29_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_29_net), 
        .M_AWADDR_28(
        PCIE_1_M_AWADDR_28_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_28_net), 
        .M_AWADDR_0(
        PCIE_1_M_AWADDR_0_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_0_net), 
        .M_AWADDR_1(
        PCIE_1_M_AWADDR_1_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_1_net), 
        .M_AWADDR_2(
        PCIE_1_M_AWADDR_2_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_2_net), 
        .M_AWADDR_3(
        PCIE_1_M_AWADDR_3_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_3_net), 
        .M_AWADDR_4(
        PCIE_1_M_AWADDR_4_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_4_net), 
        .M_AWADDR_5(
        PCIE_1_M_AWADDR_5_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_5_net), 
        .M_AWADDR_6(
        PCIE_1_M_AWADDR_6_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_6_net), 
        .M_AWADDR_7(
        PCIE_1_M_AWADDR_7_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_7_net), 
        .M_AWADDR_8(
        PCIE_1_M_AWADDR_8_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_8_net), 
        .M_AWADDR_9(
        PCIE_1_M_AWADDR_9_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_9_net), 
        .M_AWADDR_10(
        PCIE_1_M_AWADDR_10_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_10_net), 
        .M_AWADDR_11(
        PCIE_1_M_AWADDR_11_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_11_net), 
        .M_AWADDR_12(
        PCIE_1_M_AWADDR_12_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_12_net), 
        .M_AWADDR_13(
        PCIE_1_M_AWADDR_13_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_13_net), 
        .M_AWADDR_14(
        PCIE_1_M_AWADDR_14_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_14_net), 
        .M_AWADDR_15(
        PCIE_1_M_AWADDR_15_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_15_net), 
        .M_AWADDR_16(
        PCIE_1_M_AWADDR_16_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_16_net), 
        .M_AWADDR_17(
        PCIE_1_M_AWADDR_17_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_17_net), 
        .M_AWADDR_18(
        PCIE_1_M_AWADDR_18_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_18_net), 
        .M_AWADDR_19(
        PCIE_1_M_AWADDR_19_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_19_net), 
        .M_AWADDR_20(
        PCIE_1_M_AWADDR_20_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_20_net), 
        .M_AWADDR_21(
        PCIE_1_M_AWADDR_21_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_21_net), 
        .M_AWADDR_22(
        PCIE_1_M_AWADDR_22_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_22_net), 
        .M_AWADDR_23(
        PCIE_1_M_AWADDR_23_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_23_net), 
        .M_RDATA({
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_63, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_62, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_61, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_60, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_59, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_58, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_57, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_56, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_55, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_54, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_53, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_52, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_51, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_50, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_49, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_48, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_47, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_46, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_45, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_44, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_43, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_42, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_41, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_40, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_39, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_38, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_37, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_36, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_35, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_34, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_33, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_32, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_31, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_30, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_29, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_28, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_27, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_26, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_25, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_24, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_23, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_22, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_21, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_20, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_19, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_18, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_17, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_16, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_15, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_14, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_13, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_12, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_11, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_10, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_9, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_8, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_7, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_6, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_5, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_4, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_3, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_2, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_1, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_0}), 
        .M_WDATA({
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_63, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_62, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_61, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_60, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_59, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_58, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_57, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_56, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_55, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_54, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_53, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_52, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_51, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_50, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_49, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_48, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_47, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_46, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_45, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_44, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_43, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_42, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_41, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_40, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_39, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_38, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_37, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_36, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_35, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_34, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_33, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_32, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_31, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_30, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_29, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_28, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_27, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_26, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_25, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_24, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_23, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_22, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_21, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_20, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_19, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_18, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_17, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_16, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_15, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_14, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_13, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_12, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_11, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_10, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_9, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_8, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_7, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_6, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_5, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_4, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_3, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_2, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_1, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_0}), 
        .S_ARADDR_31(
        PCIE_1_S_ARADDR_31_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_31_net), 
        .S_ARADDR_30(
        PCIE_1_S_ARADDR_30_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_30_net), 
        .S_ARADDR_28(
        PCIE_1_S_ARADDR_28_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_28_net), 
        .S_ARADDR_0(
        PCIE_1_S_ARADDR_0_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_0_net), 
        .S_ARADDR_1(
        PCIE_1_S_ARADDR_1_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_1_net), 
        .S_ARADDR_2(
        PCIE_1_S_ARADDR_2_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_2_net), 
        .S_ARADDR_3(
        PCIE_1_S_ARADDR_3_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_3_net), 
        .S_ARADDR_4(
        PCIE_1_S_ARADDR_4_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_4_net), 
        .S_ARADDR_5(
        PCIE_1_S_ARADDR_5_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_5_net), 
        .S_ARADDR_6(
        PCIE_1_S_ARADDR_6_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_6_net), 
        .S_ARADDR_7(
        PCIE_1_S_ARADDR_7_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_7_net), 
        .S_ARADDR_8(
        PCIE_1_S_ARADDR_8_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_8_net), 
        .S_ARADDR_9(
        PCIE_1_S_ARADDR_9_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_9_net), 
        .S_ARADDR_10(
        PCIE_1_S_ARADDR_10_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_10_net), 
        .S_ARADDR_11(
        PCIE_1_S_ARADDR_11_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_11_net), 
        .S_ARADDR_12(
        PCIE_1_S_ARADDR_12_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_12_net), 
        .S_ARADDR_13(
        PCIE_1_S_ARADDR_13_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_13_net), 
        .S_ARADDR_14(
        PCIE_1_S_ARADDR_14_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_14_net), 
        .S_ARADDR_15(
        PCIE_1_S_ARADDR_15_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_15_net), 
        .S_ARADDR_16(
        PCIE_1_S_ARADDR_16_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_16_net), 
        .S_ARADDR_17(
        PCIE_1_S_ARADDR_17_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_17_net), 
        .S_ARADDR_18(
        PCIE_1_S_ARADDR_18_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_18_net), 
        .S_ARADDR_19(
        PCIE_1_S_ARADDR_19_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_19_net), 
        .S_ARADDR_20(
        PCIE_1_S_ARADDR_20_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_20_net), 
        .S_ARADDR_21(
        PCIE_1_S_ARADDR_21_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_21_net), 
        .S_ARADDR_22(
        PCIE_1_S_ARADDR_22_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_22_net), 
        .S_ARADDR_23(
        PCIE_1_S_ARADDR_23_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_23_net), 
        .S_AWADDR_31(
        PCIE_1_S_AWADDR_31_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_31_net), 
        .S_AWADDR_30(
        PCIE_1_S_AWADDR_30_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_30_net), 
        .S_AWADDR_28(
        PCIE_1_S_AWADDR_28_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_28_net), 
        .S_AWADDR_0(
        PCIE_1_S_AWADDR_0_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_0_net), 
        .S_AWADDR_1(
        PCIE_1_S_AWADDR_1_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_1_net), 
        .S_AWADDR_2(
        PCIE_1_S_AWADDR_2_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_2_net), 
        .S_AWADDR_3(
        PCIE_1_S_AWADDR_3_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_3_net), 
        .S_AWADDR_4(
        PCIE_1_S_AWADDR_4_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_4_net), 
        .S_AWADDR_5(
        PCIE_1_S_AWADDR_5_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_5_net), 
        .S_AWADDR_6(
        PCIE_1_S_AWADDR_6_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_6_net), 
        .S_AWADDR_7(
        PCIE_1_S_AWADDR_7_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_7_net), 
        .S_AWADDR_8(
        PCIE_1_S_AWADDR_8_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_8_net), 
        .S_AWADDR_9(
        PCIE_1_S_AWADDR_9_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_9_net), 
        .S_AWADDR_10(
        PCIE_1_S_AWADDR_10_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_10_net), 
        .S_AWADDR_11(
        PCIE_1_S_AWADDR_11_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_11_net), 
        .S_AWADDR_12(
        PCIE_1_S_AWADDR_12_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_12_net), 
        .S_AWADDR_13(
        PCIE_1_S_AWADDR_13_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_13_net), 
        .S_AWADDR_14(
        PCIE_1_S_AWADDR_14_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_14_net), 
        .S_AWADDR_15(
        PCIE_1_S_AWADDR_15_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_15_net), 
        .S_AWADDR_16(
        PCIE_1_S_AWADDR_16_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_16_net), 
        .S_AWADDR_17(
        PCIE_1_S_AWADDR_17_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_17_net), 
        .S_AWADDR_18(
        PCIE_1_S_AWADDR_18_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_18_net), 
        .S_AWADDR_19(
        PCIE_1_S_AWADDR_19_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_19_net), 
        .S_AWADDR_20(
        PCIE_1_S_AWADDR_20_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_20_net), 
        .S_AWADDR_21(
        PCIE_1_S_AWADDR_21_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_21_net), 
        .S_AWADDR_22(
        PCIE_1_S_AWADDR_22_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_22_net), 
        .S_AWADDR_23(
        PCIE_1_S_AWADDR_23_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_23_net), 
        .AXI_CLK_STABLE(AXI_CLK_STABLE_FROM_PCIECOMMON_TO_PCIE_1_net), 
        .S_RDATA({
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_63, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_62, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_61, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_60, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_59, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_58, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_57, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_56, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_55, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_54, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_53, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_52, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_51, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_50, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_49, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_48, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_47, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_46, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_45, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_44, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_43, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_42, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_41, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_40, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_39, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_38, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_37, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_36, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_35, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_34, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_33, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_32, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_31, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_30, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_29, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_28, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_27, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_26, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_25, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_24, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_23, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_22, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_21, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_20, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_19, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_18, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_17, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_16, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_15, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_14, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_13, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_12, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_11, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_10, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_9, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_8, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_7, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_6, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_5, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_4, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_3, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_2, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_1, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_0}), 
        .S_WDATA({
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_63, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_62, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_61, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_60, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_59, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_58, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_57, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_56, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_55, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_54, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_53, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_52, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_51, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_50, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_49, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_48, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_47, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_46, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_45, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_44, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_43, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_42, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_41, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_40, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_39, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_38, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_37, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_36, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_35, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_34, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_33, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_32, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_31, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_30, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_29, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_28, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_27, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_26, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_25, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_24, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_23, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_22, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_21, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_20, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_19, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_18, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_17, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_16, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_15, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_14, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_13, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_12, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_11, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_10, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_9, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_8, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_7, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_6, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_5, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_4, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_3, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_2, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_1, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_0}), 
        .PCIE_DEBUG({
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_31, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_30, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_29, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_28, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_27, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_26, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_25, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_24, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_23, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_22, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_21, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_20, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_19, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_18, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_17, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_16, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_15, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_14, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_13, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_12, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_11, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_10, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_9, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_8, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_7, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_6, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_5, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_4, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_3, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_2, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_1, 
        PCIE_1_PCIE_DEBUG_PCIE_COMMON_INSTANCE_PCIE_DEBUG_1_net_0}), 
        .DRI_CLK(), .DRI_CTRL({nc66, nc67, nc68, nc69, nc70, nc71, 
        nc72, nc73, nc74, nc75, nc76}), .DRI_WDATA({nc77, nc78, nc79, 
        nc80, nc81, nc82, nc83, nc84, nc85, nc86, nc87, nc88, nc89, 
        nc90, nc91, nc92, nc93, nc94, nc95, nc96, nc97, nc98, nc99, 
        nc100, nc101, nc102, nc103, nc104, nc105, nc106, nc107, nc108, 
        nc109}), .DRI_ARST_N(), .DRI_RDATA({nc110, nc111, nc112, nc113, 
        nc114, nc115, nc116, nc117, nc118, nc119, nc120, nc121, nc122, 
        nc123, nc124, nc125, nc126, nc127, nc128, nc129, nc130, nc131, 
        nc132, nc133, nc134, nc135, nc136, nc137, nc138, nc139, nc140, 
        nc141, nc142}), .DRI_INTERRUPT(), .DRI_BRIDGE_CLK(), 
        .DRI_BRIDGE_CTRL({nc143, nc144, nc145, nc146, nc147, nc148, 
        nc149, nc150, nc151, nc152, nc153}), .DRI_BRIDGE_WDATA({nc154, 
        nc155, nc156, nc157, nc158, nc159, nc160, nc161, nc162, nc163, 
        nc164, nc165, nc166, nc167, nc168, nc169, nc170, nc171, nc172, 
        nc173, nc174, nc175, nc176, nc177, nc178, nc179, nc180, nc181, 
        nc182, nc183, nc184, nc185, nc186}), .DRI_BRIDGE_ARST_N(), 
        .DRI_BRIDGE_RDATA({nc187, nc188, nc189, nc190, nc191, nc192, 
        nc193, nc194, nc195, nc196, nc197, nc198, nc199, nc200, nc201, 
        nc202, nc203, nc204, nc205, nc206, nc207, nc208, nc209, nc210, 
        nc211, nc212, nc213, nc214, nc215, nc216, nc217, nc218, nc219})
        , .DRI_BRIDGE_INTERRUPT(), .ARST_N({nc220, nc221, nc222, nc223})
        , .XCVR_ARST_N({vcc_net, vcc_net}), .PHYSTATUS_0(vcc_net), 
        .PHYSTATUS_1(vcc_net), .PHYSTATUS_2(
        PCIE_1_PHYSTATUS_2_PCIESS_LANE2_Pipe_AXI1_PHYSTATUS_0_net), 
        .PHYSTATUS_3(
        PCIE_1_PHYSTATUS_3_PCIESS_LANE3_Pipe_AXI0_PHYSTATUS_0_net), 
        .POWERDOWN({
        PCIE_1_POWERDOWN_PCIESS_LANE2_Pipe_AXI1_POWERDOWN_net_1, 
        PCIE_1_POWERDOWN_PCIESS_LANE2_Pipe_AXI1_POWERDOWN_net_0}), 
        .RATE({PCIE_1_RATE_PCIESS_LANE2_Pipe_AXI1_RATE_net_1, 
        PCIE_1_RATE_PCIESS_LANE2_Pipe_AXI1_RATE_net_0}), .RESET_N(
        PCIE_1_RESET_N_PCIESS_LANE2_Pipe_AXI1_RESET_N_net), .RXDATA_0({
        gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, 
        gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, 
        gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, 
        gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, 
        gnd_net, gnd_net, gnd_net, gnd_net}), .RXDATA_1({gnd_net, 
        gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, 
        gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, 
        gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, 
        gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, 
        gnd_net, gnd_net, gnd_net}), .RXDATA_2({
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_31, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_30, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_29, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_28, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_27, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_26, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_25, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_24, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_23, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_22, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_21, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_20, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_19, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_18, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_17, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_16, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_15, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_14, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_13, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_12, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_11, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_10, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_9, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_8, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_7, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_6, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_5, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_4, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_3, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_2, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_1, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_0}), 
        .RXDATA_3({
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_31, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_30, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_29, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_28, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_27, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_26, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_25, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_24, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_23, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_22, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_21, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_20, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_19, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_18, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_17, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_16, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_15, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_14, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_13, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_12, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_11, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_10, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_9, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_8, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_7, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_6, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_5, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_4, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_3, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_2, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_1, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_0}), 
        .RXDATAK_0({gnd_net, gnd_net, gnd_net, gnd_net}), .RXDATAK_1({
        gnd_net, gnd_net, gnd_net, gnd_net}), .RXDATAK_2({
        PCIE_1_RXDATAK_2_PCIESS_LANE2_Pipe_AXI1_RXDATAK_0_net_3, 
        PCIE_1_RXDATAK_2_PCIESS_LANE2_Pipe_AXI1_RXDATAK_0_net_2, 
        PCIE_1_RXDATAK_2_PCIESS_LANE2_Pipe_AXI1_RXDATAK_0_net_1, 
        PCIE_1_RXDATAK_2_PCIESS_LANE2_Pipe_AXI1_RXDATAK_0_net_0}), 
        .RXDATAK_3({
        PCIE_1_RXDATAK_3_PCIESS_LANE3_Pipe_AXI0_RXDATAK_0_net_3, 
        PCIE_1_RXDATAK_3_PCIESS_LANE3_Pipe_AXI0_RXDATAK_0_net_2, 
        PCIE_1_RXDATAK_3_PCIESS_LANE3_Pipe_AXI0_RXDATAK_0_net_1, 
        PCIE_1_RXDATAK_3_PCIESS_LANE3_Pipe_AXI0_RXDATAK_0_net_0}), 
        .RXELECIDLE_0(vcc_net), .RXELECIDLE_1(vcc_net), .RXELECIDLE_2(
        PCIE_1_RXELECIDLE_2_PCIESS_LANE2_Pipe_AXI1_RXELECIDLE_0_net), 
        .RXELECIDLE_3(
        PCIE_1_RXELECIDLE_3_PCIESS_LANE3_Pipe_AXI0_RXELECIDLE_0_net), 
        .RXPOLARITY_0(), .RXPOLARITY_1(), .RXPOLARITY_2(
        PCIE_1_RXPOLARITY_2_PCIESS_LANE2_Pipe_AXI1_RXPOLARITY_0_net), 
        .RXPOLARITY_3(
        PCIE_1_RXPOLARITY_3_PCIESS_LANE3_Pipe_AXI0_RXPOLARITY_0_net), 
        .RXSTANDBYSTATUS_0(), .RXSTANDBYSTATUS_1(), .RXSTANDBYSTATUS_2(
        PCIE_1_RXSTANDBYSTATUS_2_PCIESS_LANE2_Pipe_AXI1_RXSTANDBYSTATUS_0_net)
        , .RXSTANDBYSTATUS_3(
        PCIE_1_RXSTANDBYSTATUS_3_PCIESS_LANE3_Pipe_AXI0_RXSTANDBYSTATUS_0_net)
        , .RXSTATUS_0({gnd_net, gnd_net, gnd_net}), .RXSTATUS_1({
        gnd_net, gnd_net, gnd_net}), .RXSTATUS_2({
        PCIE_1_RXSTATUS_2_PCIESS_LANE2_Pipe_AXI1_RXSTATUS_0_net_2, 
        PCIE_1_RXSTATUS_2_PCIESS_LANE2_Pipe_AXI1_RXSTATUS_0_net_1, 
        PCIE_1_RXSTATUS_2_PCIESS_LANE2_Pipe_AXI1_RXSTATUS_0_net_0}), 
        .RXSTATUS_3({
        PCIE_1_RXSTATUS_3_PCIESS_LANE3_Pipe_AXI0_RXSTATUS_0_net_2, 
        PCIE_1_RXSTATUS_3_PCIESS_LANE3_Pipe_AXI0_RXSTATUS_0_net_1, 
        PCIE_1_RXSTATUS_3_PCIESS_LANE3_Pipe_AXI0_RXSTATUS_0_net_0}), 
        .RXVALID_0(gnd_net), .RXVALID_1(gnd_net), .RXVALID_2(
        PCIE_1_RXVALID_2_PCIESS_LANE2_Pipe_AXI1_RXVALID_0_net), 
        .RXVALID_3(
        PCIE_1_RXVALID_3_PCIESS_LANE3_Pipe_AXI0_RXVALID_0_net), 
        .TXCOMPLIANCE_0(), .TXCOMPLIANCE_1(), .TXCOMPLIANCE_2(
        PCIE_1_TXCOMPLIANCE_2_PCIESS_LANE2_Pipe_AXI1_TXCOMPLIANCE_0_net)
        , .TXCOMPLIANCE_3(
        PCIE_1_TXCOMPLIANCE_3_PCIESS_LANE3_Pipe_AXI0_TXCOMPLIANCE_0_net)
        , .TXDATA_0({nc224, nc225, nc226, nc227, nc228, nc229, nc230, 
        nc231, nc232, nc233, nc234, nc235, nc236, nc237, nc238, nc239, 
        nc240, nc241, nc242, nc243, nc244, nc245, nc246, nc247, nc248, 
        nc249, nc250, nc251, nc252, nc253, nc254, nc255}), .TXDATA_1({
        nc256, nc257, nc258, nc259, nc260, nc261, nc262, nc263, nc264, 
        nc265, nc266, nc267, nc268, nc269, nc270, nc271, nc272, nc273, 
        nc274, nc275, nc276, nc277, nc278, nc279, nc280, nc281, nc282, 
        nc283, nc284, nc285, nc286, nc287}), .TXDATA_2({
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_31, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_30, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_29, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_28, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_27, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_26, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_25, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_24, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_23, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_22, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_21, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_20, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_19, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_18, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_17, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_16, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_15, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_14, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_13, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_12, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_11, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_10, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_9, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_8, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_7, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_6, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_5, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_4, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_3, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_2, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_1, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_0}), 
        .TXDATA_3({
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_31, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_30, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_29, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_28, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_27, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_26, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_25, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_24, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_23, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_22, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_21, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_20, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_19, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_18, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_17, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_16, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_15, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_14, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_13, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_12, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_11, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_10, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_9, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_8, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_7, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_6, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_5, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_4, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_3, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_2, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_1, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_0}), 
        .TXDATAK_0({nc288, nc289, nc290, nc291}), .TXDATAK_1({nc292, 
        nc293, nc294, nc295}), .TXDATAK_2({
        PCIE_1_TXDATAK_2_PCIESS_LANE2_Pipe_AXI1_TXDATAK_0_net_3, 
        PCIE_1_TXDATAK_2_PCIESS_LANE2_Pipe_AXI1_TXDATAK_0_net_2, 
        PCIE_1_TXDATAK_2_PCIESS_LANE2_Pipe_AXI1_TXDATAK_0_net_1, 
        PCIE_1_TXDATAK_2_PCIESS_LANE2_Pipe_AXI1_TXDATAK_0_net_0}), 
        .TXDATAK_3({
        PCIE_1_TXDATAK_3_PCIESS_LANE3_Pipe_AXI0_TXDATAK_0_net_3, 
        PCIE_1_TXDATAK_3_PCIESS_LANE3_Pipe_AXI0_TXDATAK_0_net_2, 
        PCIE_1_TXDATAK_3_PCIESS_LANE3_Pipe_AXI0_TXDATAK_0_net_1, 
        PCIE_1_TXDATAK_3_PCIESS_LANE3_Pipe_AXI0_TXDATAK_0_net_0}), 
        .TXDATAVALID_0(), .TXDATAVALID_1(), .TXDATAVALID_2(
        PCIE_1_TXDATAVALID_2_PCIESS_LANE2_Pipe_AXI1_TXDATAVALID_0_net), 
        .TXDATAVALID_3(
        PCIE_1_TXDATAVALID_3_PCIESS_LANE3_Pipe_AXI0_TXDATAVALID_0_net), 
        .TXDEEMPH(PCIE_1_TXDEEMPH_PCIESS_LANE2_Pipe_AXI1_TXDEEMPH_net), 
        .TXDETECTRX_LOOPBACK_0(), .TXDETECTRX_LOOPBACK_1(), 
        .TXDETECTRX_LOOPBACK_2(
        PCIE_1_TXDETECTRX_LOOPBACK_2_PCIESS_LANE2_Pipe_AXI1_TXDETECTRX_LOOPBACK_0_net)
        , .TXDETECTRX_LOOPBACK_3(
        PCIE_1_TXDETECTRX_LOOPBACK_3_PCIESS_LANE3_Pipe_AXI0_TXDETECTRX_LOOPBACK_0_net)
        , .TXELECIDLE_0(), .TXELECIDLE_1(), .TXELECIDLE_2(
        PCIE_1_TXELECIDLE_2_PCIESS_LANE2_Pipe_AXI1_TXELECIDLE_0_net), 
        .TXELECIDLE_3(
        PCIE_1_TXELECIDLE_3_PCIESS_LANE3_Pipe_AXI0_TXELECIDLE_0_net), 
        .TXMARGIN({
        PCIE_1_TXMARGIN_PCIESS_LANE2_Pipe_AXI1_TXMARGIN_net_2, 
        PCIE_1_TXMARGIN_PCIESS_LANE2_Pipe_AXI1_TXMARGIN_net_1, 
        PCIE_1_TXMARGIN_PCIESS_LANE2_Pipe_AXI1_TXMARGIN_net_0}), 
        .TXSWING(PCIE_1_TXSWING_PCIESS_LANE2_Pipe_AXI1_TXSWING_net), 
        .PIPE_CLK_0(), .PIPE_CLK_1(), .PIPE_CLK_2(
        PCIE_1_PIPE_CLK_2_PCIESS_LANE2_Pipe_AXI1_PIPE_CLK_0_net), 
        .PIPE_CLK_3(
        PCIE_1_PIPE_CLK_3_PCIESS_LANE3_Pipe_AXI0_PIPE_CLK_0_net), 
        .PCLK_OUT_0(gnd_net), .PCLK_OUT_1(gnd_net), .PCLK_OUT_2(
        PCIE_1_PCLK_OUT_2_PCIESS_LANE2_Pipe_AXI1_PCLK_OUT_0_net), 
        .PCLK_OUT_3(
        PCIE_1_PCLK_OUT_3_PCIESS_LANE3_Pipe_AXI0_PCLK_OUT_0_net), 
        .AXI_CLK(PCIE_COMMON_AXI_CLK_OUT_net), .LINK_BRIDGE_CLK(
        pcie_apblink_inst_PCIE1_BRIDGE_CLK_PCIE_1_LINK_BRIDGE_CLK_net), 
        .LINK_BRIDGE_ADDR({
        pcie_apblink_inst_PCIE1_BRIDGE_ADDR_PCIE_1_LINK_BRIDGE_ADDR_net_2, 
        pcie_apblink_inst_PCIE1_BRIDGE_ADDR_PCIE_1_LINK_BRIDGE_ADDR_net_1, 
        pcie_apblink_inst_PCIE1_BRIDGE_ADDR_PCIE_1_LINK_BRIDGE_ADDR_net_0})
        , .LINK_BRIDGE_EN(
        pcie_apblink_inst_PCIE1_BRIDGE_EN_PCIE_1_LINK_BRIDGE_EN_net), 
        .LINK_BRIDGE_ARST_N(
        pcie_apblink_inst_PCIE1_BRIDGE_ARST_N_PCIE_1_LINK_BRIDGE_ARST_N_net)
        , .LINK_BRIDGE_WDATA({
        pcie_apblink_inst_PCIE1_BRIDGE_WDATA_PCIE_1_LINK_BRIDGE_WDATA_net_3, 
        pcie_apblink_inst_PCIE1_BRIDGE_WDATA_PCIE_1_LINK_BRIDGE_WDATA_net_2, 
        pcie_apblink_inst_PCIE1_BRIDGE_WDATA_PCIE_1_LINK_BRIDGE_WDATA_net_1, 
        pcie_apblink_inst_PCIE1_BRIDGE_WDATA_PCIE_1_LINK_BRIDGE_WDATA_net_0})
        , .LINK_BRIDGE_RDATA({
        pcie_apblink_inst_PCIE1_BRIDGE_RDATA_PCIE_1_LINK_BRIDGE_RDATA_net_3, 
        pcie_apblink_inst_PCIE1_BRIDGE_RDATA_PCIE_1_LINK_BRIDGE_RDATA_net_2, 
        pcie_apblink_inst_PCIE1_BRIDGE_RDATA_PCIE_1_LINK_BRIDGE_RDATA_net_1, 
        pcie_apblink_inst_PCIE1_BRIDGE_RDATA_PCIE_1_LINK_BRIDGE_RDATA_net_0})
        , .LINK_CTRL_CLK(gnd_net), .LINK_CTRL_ADDR({gnd_net, gnd_net, 
        gnd_net}), .LINK_CTRL_EN(gnd_net), .LINK_CTRL_ARST_N(gnd_net), 
        .LINK_CTRL_WDATA({gnd_net, gnd_net, gnd_net, gnd_net}), 
        .LINK_CTRL_RDATA({nc296, nc297, nc298, nc299}));
    G5_APBLINK_MASTER pcie_apblink_master_inst (.preset_b(
        APB_S_PRESET_N), .pclk(APB_S_PCLK), .psel(APB_S_PSEL), 
        .penable(APB_S_PENABLE), .pwrite(APB_S_PWRITE), .pstrb({
        vcc_net, vcc_net, vcc_net, vcc_net}), .paddr({APB_S_PADDR[27], 
        APB_S_PADDR[26], APB_S_PADDR[25], APB_S_PADDR[24], 
        APB_S_PADDR[23], APB_S_PADDR[22], APB_S_PADDR[21], 
        APB_S_PADDR[20], APB_S_PADDR[19], APB_S_PADDR[18], 
        APB_S_PADDR[17], APB_S_PADDR[16], APB_S_PADDR[15], 
        APB_S_PADDR[14], APB_S_PADDR[13], APB_S_PADDR[12], 
        APB_S_PADDR[11], APB_S_PADDR[10], APB_S_PADDR[9], 
        APB_S_PADDR[8], APB_S_PADDR[7], APB_S_PADDR[6], APB_S_PADDR[5], 
        APB_S_PADDR[4], APB_S_PADDR[3], APB_S_PADDR[2]}), .pwdata({
        APB_S_PWDATA[31], APB_S_PWDATA[30], APB_S_PWDATA[29], 
        APB_S_PWDATA[28], APB_S_PWDATA[27], APB_S_PWDATA[26], 
        APB_S_PWDATA[25], APB_S_PWDATA[24], APB_S_PWDATA[23], 
        APB_S_PWDATA[22], APB_S_PWDATA[21], APB_S_PWDATA[20], 
        APB_S_PWDATA[19], APB_S_PWDATA[18], APB_S_PWDATA[17], 
        APB_S_PWDATA[16], APB_S_PWDATA[15], APB_S_PWDATA[14], 
        APB_S_PWDATA[13], APB_S_PWDATA[12], APB_S_PWDATA[11], 
        APB_S_PWDATA[10], APB_S_PWDATA[9], APB_S_PWDATA[8], 
        APB_S_PWDATA[7], APB_S_PWDATA[6], APB_S_PWDATA[5], 
        APB_S_PWDATA[4], APB_S_PWDATA[3], APB_S_PWDATA[2], 
        APB_S_PWDATA[1], APB_S_PWDATA[0]}), .lnk_m_rdata({
        pcie_apblink_master_inst_lnk_m_rdata_pcie_apblink_inst_S_RDATA_net_3, 
        pcie_apblink_master_inst_lnk_m_rdata_pcie_apblink_inst_S_RDATA_net_2, 
        pcie_apblink_master_inst_lnk_m_rdata_pcie_apblink_inst_S_RDATA_net_1, 
        pcie_apblink_master_inst_lnk_m_rdata_pcie_apblink_inst_S_RDATA_net_0})
        , .pready(APB_S_PREADY), .pslverr(APB_S_PSLVERR), .lnk_m_rst_b(
        pcie_apblink_master_inst_lnk_m_rst_b_pcie_apblink_inst_S_ARST_N_net)
        , .lnk_m_enable(
        pcie_apblink_master_inst_lnk_m_enable_pcie_apblink_inst_S_EN_net)
        , .lnk_m_clock(
        pcie_apblink_master_inst_lnk_m_clock_pcie_apblink_inst_S_CLK_net)
        , .lnk_m_addr({
        pcie_apblink_master_inst_lnk_m_addr_pcie_apblink_inst_S_ADDR_net_2, 
        pcie_apblink_master_inst_lnk_m_addr_pcie_apblink_inst_S_ADDR_net_1, 
        pcie_apblink_master_inst_lnk_m_addr_pcie_apblink_inst_S_ADDR_net_0})
        , .lnk_m_wdata({
        pcie_apblink_master_inst_lnk_m_wdata_pcie_apblink_inst_S_WDATA_net_3, 
        pcie_apblink_master_inst_lnk_m_wdata_pcie_apblink_inst_S_WDATA_net_2, 
        pcie_apblink_master_inst_lnk_m_wdata_pcie_apblink_inst_S_WDATA_net_1, 
        pcie_apblink_master_inst_lnk_m_wdata_pcie_apblink_inst_S_WDATA_net_0})
        , .lnk_state_copy({nc300, nc301, nc302, nc303, nc304, nc305}), 
        .prdata({APB_S_PRDATA[31], APB_S_PRDATA[30], APB_S_PRDATA[29], 
        APB_S_PRDATA[28], APB_S_PRDATA[27], APB_S_PRDATA[26], 
        APB_S_PRDATA[25], APB_S_PRDATA[24], APB_S_PRDATA[23], 
        APB_S_PRDATA[22], APB_S_PRDATA[21], APB_S_PRDATA[20], 
        APB_S_PRDATA[19], APB_S_PRDATA[18], APB_S_PRDATA[17], 
        APB_S_PRDATA[16], APB_S_PRDATA[15], APB_S_PRDATA[14], 
        APB_S_PRDATA[13], APB_S_PRDATA[12], APB_S_PRDATA[11], 
        APB_S_PRDATA[10], APB_S_PRDATA[9], APB_S_PRDATA[8], 
        APB_S_PRDATA[7], APB_S_PRDATA[6], APB_S_PRDATA[5], 
        APB_S_PRDATA[4], APB_S_PRDATA[3], APB_S_PRDATA[2], 
        APB_S_PRDATA[1], APB_S_PRDATA[0]}));
    GND PCIESS_AXI_1_M_AWLEN_5_GndInst (.Y(PCIESS_AXI_1_M_AWLEN[5]));
    XCVR_PIPE_AXI0 #( .MAIN_QMUX_R0_QRST0_SRC(3'b001), .MAIN_QMUX_R0_QRST1_SRC(3'b011)
        , .MAIN_QMUX_R0_QRST2_SRC(3'b000), .MAIN_QMUX_R0_QRST3_SRC(3'b000)
        , .DATA_RATE(5000.0), .REG_FILE(""), .PMA_CMN_SOFT_RESET_NV_MAP(1'b0)
        , .PMA_CMN_SOFT_RESET_V_MAP(1'b0), .PMA_CMN_SOFT_RESET_PERIPH(1'b0)
        , .PMA_CMN_TXPLL_CLKBUF_TXPLL_DUALCLK1_MODE(2'b00), .PMA_CMN_TXPLL_CLKBUF_TXPLL_DUALCLK1_ENTERM(2'b00)
        , .PMA_CMN_TXPLL_CLKBUF_TXPLL_DUALCLK0_MODE(2'b10), .PMA_CMN_TXPLL_CLKBUF_TXPLL_DUALCLK0_ENTERM(2'b00)
        , .PMA_CMN_TXPLL_CLKBUF_TXPLL_DUALCLK1_EN_HYST(1'b0), .PMA_CMN_TXPLL_CLKBUF_TXPLL_DUALCLK0_EN_HYST(1'b0)
        , .PMA_CMN_TXPLL_CLKBUF_TXPLL_CLKBUF_EN_RDIFF(1'b0), .PMA_CMN_TXPLL_CLKBUF_TXPLL_CLKBUF_EN_UDRIVE_P(1'b1)
        , .PMA_CMN_TXPLL_CLKBUF_TXPLL_CLKBUF_EN_UDRIVE_N(1'b1), .PMA_CMN_TXPLL_CLKBUF_TXPLL_CLKBUF_EN_PULLUP(1'b0)
        , .PMA_CMN_TXPLL_CLKBUF_TXPLL_CLKBUF_EN_APAD(1'b0), .PMA_CMN_TXPLL_CTRL_TXPLL_BWSEL(1'b1)
        , .PMA_CMN_TXPLL_CTRL_TXPLL_VBGREF_SEL(1'b0), .PMA_CMN_TXPLL_CTRL_TXPLL_FBDIV_SEL(2'b00)
        , .PMA_CMN_TXPLL_CTRL_TXPLL_DSMPD(1'b0), .PMA_CMN_TXPLL_CTRL_TXPLL_PHASESTEPAMOUNT(8'b00000110)
        , .PMA_CMN_TXPLL_CTRL_TXPLL_STEP_PHASE(1'b0), .PMA_CMN_TXPLL_CTRL_TXPLL_PD(1'b0)
        , .PMA_CMN_TXPLL_CTRL_TXPLL_AUXDIVPD(1'b0), .PMA_CMN_TXPLL_CTRL_TXPLL_CLKRESETEN(1'b0)
        , .PMA_CMN_TXPLL_CTRL_TXPLL_CLKRESET(1'b0), .PMA_CMN_TXPLL_CTRL_RESET_RTL_TXPLL(1'b0)
        , .PMA_CMN_TXPLL_CTRL_RESET_RTL(1'b0), .PMA_CMN_TXPLL_CTRL_TXPLL_FOUTAUXDIV2_SEL(1'b0)
        , .PMA_CMN_TXPLL_CLK_SEL_TXPLL_REFCLK_SEL_HM(2'b11), .PMA_CMN_TXPLL_CLK_SEL_TXPLL_REFCLK_SEL_SM(3'b000)
        , .PMA_CMN_TXPLL_CLK_SEL_CASCADE_CLK_SEL_HM(2'b00), .PMA_CMN_TXPLL_CLK_SEL_CASCADE_CLK_SEL_SM(3'b111)
        , .PMA_CMN_TXPLL_CLK_SEL_TXPLL_JA_FREF_SEL(3'b000), .PMA_CMN_TXPLL_CLK_SEL_CDRCLK_LN01_INT_SEL(3'b111)
        , .PMA_CMN_TXPLL_CLK_SEL_CDRCLK_LN23_INT_SEL(3'b111), .PMA_CMN_TXPLL_CLK_SEL_CDRCLK_OUT_UP_SEL(3'b111)
        , .PMA_CMN_TXPLL_CLK_SEL_CDRCLK_OUT_DN_SEL(3'b111), .PMA_CMN_TXPLL_DIV_1_TXPLL_AUXDIV(12'b000000011001)
        , .PMA_CMN_TXPLL_DIV_1_TXPLL_FBDIV(12'b000000011001), .PMA_CMN_TXPLL_DIV_2_TXPLL_FRAC(24'b000000000000000000000001)
        , .PMA_CMN_TXPLL_DIV_2_TXPLL_REFDIV(6'b000001), .PMA_CMN_TXPLL_JA_1_TXPLL_JA_DIVFIN(16'b0000000001100100)
        , .PMA_CMN_TXPLL_JA_1_TXPLL_JA_DIVFFB(16'b0000000001100100), .PMA_CMN_TXPLL_JA_2_TXPLL_JA_SYNCCNTMAX(32'b00000000000000000000000001100100)
        , .PMA_CMN_TXPLL_JA_3_TXPLL_JA_CNTOFFSET(16'b0000000001100100)
        , .PMA_CMN_TXPLL_JA_3_TXPLL_JA_TARGETCNT(32'b00000000000000000000000001100100)
        , .PMA_CMN_TXPLL_JA_4_TXPLL_JA_OTDLY(16'b0000000000000001), .PMA_CMN_TXPLL_JA_4_TXPLL_JA_FMI(8'b00000001)
        , .PMA_CMN_TXPLL_JA_4_TXPLL_JA_FKI(4'b0001), .PMA_CMN_TXPLL_JA_5_TXPLL_JA_PMP1(8'b00000001)
        , .PMA_CMN_TXPLL_JA_5_TXPLL_JA_PMP2(8'b00000001), .PMA_CMN_TXPLL_JA_5_TXPLL_JA_PMI1(8'b00000001)
        , .PMA_CMN_TXPLL_JA_5_TXPLL_JA_PMI2(8'b00000001), .PMA_CMN_TXPLL_JA_6_TXPLL_JA_PKP1(5'b00001)
        , .PMA_CMN_TXPLL_JA_6_TXPLL_JA_PKP2(5'b00001), .PMA_CMN_TXPLL_JA_6_TXPLL_JA_PKI1(5'b00001)
        , .PMA_CMN_TXPLL_JA_6_TXPLL_JA_PKI2(5'b00001), .PMA_CMN_TXPLL_JA_7_TXPLL_JA_DELAYK(24'b000000000000000000000001)
        , .PMA_CMN_TXPLL_JA_7_TXPLL_JA_FDONLY(1'b1), .PMA_CMN_TXPLL_JA_7_TXPLL_JA_ONTARGETOV(1'b1)
        , .PMA_CMN_TXPLL_JA_7_TXPLL_JA_PROGRAM(1'b1), .PMA_CMN_TXPLL_JA_8_TXPLL_JA_FRAC_PRESET(24'b000000000000000000000000)
        , .PMA_CMN_TXPLL_JA_8_TXPLL_JA_PRESET_EN(1'b0), .PMA_CMN_TXPLL_JA_8_TXPLL_JA_HOLD(1'b0)
        , .PMA_CMN_TXPLL_JA_9_TXPLL_JA_INT_PRESET(12'b000000010100), .PMA_CMN_TXPLL_JA_RST_TXPLL_JA_RESET(1'b1)
        , .PMA_CMN_TXPLL_JA_RST_TXPLL_JA_RESET_FFB_OVERRIDE(1'b0), .PMA_CMN_TXPLL_JA_RST_TXPLL_JA_RESET_FFB_EXT(1'b1)
        , .PMA_CMN_TXPLL_JA_RST_TXPLL_JA_RESET_FIN_OVERRIDE(1'b0), .PMA_CMN_TXPLL_JA_RST_TXPLL_JA_RESET_FIN_EXT(1'b1)
        , .PMA_CMN_TXPLL_JA_RST_TXPLL_JA_RESET_CLKS_OVERRIDE(1'b0), .PMA_CMN_TXPLL_JA_RST_TXPLL_JA_RESET_CLKS_EXT(1'b1)
        , .PMA_CMN_SERDES_SSMOD_SSMOD_DOWNSPREAD(1'b0), .PMA_CMN_SERDES_SSMOD_SSMOD_DISABLE_SSCG(1'b1)
        , .PMA_CMN_SERDES_SSMOD_SSMOD_SPREAD(5'b00000), .PMA_CMN_SERDES_SSMOD_SSMOD_DIVVAL(6'b000001)
        , .PMA_CMN_SERDES_SSMOD_SSMOD_EXT_MAXADDR(8'b01111111), .PMA_CMN_SERDES_SSMOD_SSMOD_SEL_EXTWAVE(2'b00)
        , .PMA_CMN_SERDES_SSMOD_RN_SEL(2'b00), .PMA_CMN_SERDES_SSMOD_RN_FILTER(1'b0)
        , .PMA_CMN_SERDES_RTERM_RTERMCAL85(4'b0011), .PMA_CMN_SERDES_RTERM_RTERMCAL100(4'b0111)
        , .PMA_CMN_SERDES_RTERM_RTERMCAL150(4'b1101), .PMA_CMN_SERDES_RTT_RTT_CAL_TERM(4'b0000)
        , .PMA_CMN_SERDES_RTT_RTT_CURRENT_PROG(2'b00), .PMA_SOFT_RESET_NV_MAP(1'b0)
        , .PMA_SOFT_RESET_V_MAP(1'b0), .PMA_DES_CDR_CTRL_1_DCFBEN_CDR(1'b0)
        , .PMA_DES_CDR_CTRL_1_H0CDR0(5'b00000), .PMA_DES_CDR_CTRL_1_H0CDR1(5'b00000)
        , .PMA_DES_CDR_CTRL_1_H0CDR2(8'b00000000), .PMA_DES_CDR_CTRL_1_H0CDR3(5'b00000)
        , .PMA_DES_CDR_CTRL_1_CMRTRIM_CDR(3'b000), .PMA_DES_CDR_CTRL_2_CSENT1_CDR(2'b01)
        , .PMA_DES_CDR_CTRL_2_CSENT2_CDR(2'b01), .PMA_DES_CDR_CTRL_2_CSENT3_CDR(2'b01)
        , .PMA_DES_CDR_CTRL_3_SLIP_DES_CDR(1'b0), .PMA_DES_CDR_CTRL_3_SLIP_DES_CDR_SEL(1'b0)
        , .PMA_DES_CDR_CTRL_3_SLIP_DES_CDR_EN(1'b0), .PMA_DES_DFEEM_CTRL_1_CSENT1_DFEEM(2'b01)
        , .PMA_DES_DFEEM_CTRL_1_CSENT2_DFEEM(2'b01), .PMA_DES_DFEEM_CTRL_1_CSENT3_DFEEM(2'b01)
        , .PMA_DES_DFEEM_CTRL_1_CMRTRIM_DFEEM(3'b000), .PMA_DES_DFEEM_CTRL_2_H1(5'b00000)
        , .PMA_DES_DFEEM_CTRL_2_H2(5'b00000), .PMA_DES_DFEEM_CTRL_2_H3(5'b00000)
        , .PMA_DES_DFEEM_CTRL_2_H4(5'b00000), .PMA_DES_DFEEM_CTRL_3_H5(5'b00000)
        , .PMA_DES_DFE_CTRL_1_DCFBEN_DFE(1'b0), .PMA_DES_DFE_CTRL_1_H0DFE0(5'b00000)
        , .PMA_DES_DFE_CTRL_1_H0DFE1(5'b00000), .PMA_DES_DFE_CTRL_2_PHICTRL_TH_DFE(8'b00000000)
        , .PMA_DES_DFE_CTRL_2_PHICTRL_GRAY_DFE(3'b000), .PMA_DES_DFE_CTRL_2_SLIP_DES_DFE(1'b0)
        , .PMA_DES_DFE_CTRL_2_SLIP_DES_DFE_SEL(1'b0), .PMA_DES_DFE_CTRL_2_SLIP_DES_DFE_EN(1'b0)
        , .PMA_DES_EM_CTRL_1_DCFBEN_EM(1'b0), .PMA_DES_EM_CTRL_1_H0EM0(5'b00000)
        , .PMA_DES_EM_CTRL_1_H0EM1(5'b00000), .PMA_DES_EM_CTRL_1_CALIBRATION_CLK_EN(1'b0)
        , .PMA_DES_EM_CTRL_2_PHICTRL_TH_EM(8'b00000000), .PMA_DES_EM_CTRL_2_PHICTRL_GRAY_EM(3'b000)
        , .PMA_DES_EM_CTRL_2_SLIP_DES_EM(1'b0), .PMA_DES_EM_CTRL_2_SLIP_DES_EM_SEL(1'b0)
        , .PMA_DES_EM_CTRL_2_SLIP_DES_EM_EN(1'b0), .PMA_DES_RTL_EM_RUN_EYEMONITOR_COMPARISON(1'b0)
        , .PMA_DES_RTL_EM_EYEMONITOR_SAMPLE_COUNT(12'b000001100100), .PMA_DES_RTL_LOCK_CTRL_LOCK_OVERRIDE_FROMFAB(1'b0)
        , .PMA_DES_TEST_BUS_RXATESTSEL(3'b000), .PMA_DES_TEST_BUS_RXDTESTEN(1'b0)
        , .PMA_DES_TEST_BUS_RXDTESTSEL(3'b000), .PMA_DES_CLK_CTRL_RXBYPASSEN(1'b0)
        , .PMA_DES_RSTPD_RXPD(1'b0), .PMA_DES_RSTPD_RESETDES(1'b0), .PMA_DES_RSTPD_PDDFE(1'b1)
        , .PMA_DES_RSTPD_PDEM(1'b1), .PMA_DES_RSTPD_RCVEN(1'b1), .PMA_DES_RSTPD_RESET_FIFO(1'b0)
        , .PMA_DES_RTL_ERR_CHK_READ_ERROR(1'b0), .PMA_DES_PCIE1_2_RXPLL_DIV_PCIE1_RXPLL_FBDIV(8'b00011001)
        , .PMA_DES_PCIE1_2_RXPLL_DIV_PCIE1_RXPLL_REFDIV(5'b00010), .PMA_DES_PCIE1_2_RXPLL_DIV_PCIE1_RXPLL_RANGE(2'b01)
        , .PMA_DES_PCIE1_2_RXPLL_DIV_PCIE2_RXPLL_FBDIV(8'b00110010), .PMA_DES_PCIE1_2_RXPLL_DIV_PCIE2_RXPLL_REFDIV(5'b00010)
        , .PMA_DES_PCIE1_2_RXPLL_DIV_PCIE2_RXPLL_RANGE(2'b00), .PMA_DES_SATA1_2_RXPLL_DIV_SATA1_RXPLL_FBDIV(8'b00011000)
        , .PMA_DES_SATA1_2_RXPLL_DIV_SATA1_RXPLL_REFDIV(5'b00100), .PMA_DES_SATA1_2_RXPLL_DIV_SATA1_RXPLL_RANGE(2'b10)
        , .PMA_DES_SATA1_2_RXPLL_DIV_SATA2_RXPLL_FBDIV(8'b00011000), .PMA_DES_SATA1_2_RXPLL_DIV_SATA2_RXPLL_REFDIV(5'b00010)
        , .PMA_DES_SATA1_2_RXPLL_DIV_SATA2_RXPLL_RANGE(2'b01), .PMA_DES_SATA3_RXPLL_DIV_SATA3_RXPLL_FBDIV(8'b00110000)
        , .PMA_DES_SATA3_RXPLL_DIV_SATA3_RXPLL_REFDIV(5'b00010), .PMA_DES_SATA3_RXPLL_DIV_SATA3_RXPLL_RANGE(2'b00)
        , .PMA_SER_CTRL_CMSTEP_VALUE(1'b0), .PMA_SER_CTRL_CMSTEP(1'b0)
        , .PMA_SER_CTRL_NLPBK_EN(1'b0), .PMA_SER_CTRL_HSLPBKEN(1'b0), .PMA_SER_CTRL_HSLPBK_SEL(3'b000)
        , .PMA_SER_RSTPD_RESETSEREN(1'b1), .PMA_SER_RSTPD_RESETSER(1'b0)
        , .PMA_SER_RSTPD_TXPD(1'b0), .PMA_SER_DRV_BYP_BYPASSSER(1'b0)
        , .PMA_SER_RXDET_CTRL_RXDETECT_COUNT_THRESHOLD(14'b00000000000001)
        , .PMA_SER_RXDET_CTRL_RX_DETECT_EN(1'b0), .PMA_SER_RXDET_CTRL_RXDETECT_START(1'b0)
        , .PMA_SER_STATIC_LSB_STATIC_PATTERN_LSB(20'b00000000000000000000)
        , .PMA_SER_STATIC_MSB_STATIC_PATTERN_MSB(20'b00000000000000000000)
        , .PMA_SER_TEST_BUS_TXATESTSEL(3'b000), .PMA_SER_TEST_BUS_DTESTEN_RTL(1'b0)
        , .PMA_SER_TEST_BUS_DTESTSEL_RTL(4'b0000), .PMA_SER_TEST_BUS_JTAG_TO_DTEST_SEL(3'b000)
        , .PMA_SER_TEST_BUS_PRBSERR_TO_DTEST_SEL(2'b00), .PMA_SER_TEST_BUS_RXPKDETOUT_TO_DTEST_SEL(3'b111)
        , .PMA_SER_DRV_CTRL_M0_TXDRVTRIM_FS_3P5DB_M0(6'b100011), .PMA_SER_DRV_CTRL_M0_TXDRVTRIM_FS_6P0DB_M0(6'b110100)
        , .PMA_SER_DRV_CTRL_M0_TXDRVTRIM_HS_0DB_M0(6'b011011), .PMA_SER_DRV_CTRL_M1_TXDRVTRIM_FS_3P5DB_M1(6'b100111)
        , .PMA_SER_DRV_CTRL_M1_TXDRVTRIM_FS_6P0DB_M1(6'b101100), .PMA_SER_DRV_CTRL_M1_TXDRVTRIM_HS_0DB_M1(6'b100011)
        , .PMA_SER_DRV_CTRL_M2_TXDRVTRIM_FS_3P5DB_M2(6'b011011), .PMA_SER_DRV_CTRL_M2_TXDRVTRIM_FS_6P0DB_M2(6'b011011)
        , .PMA_SER_DRV_CTRL_M2_TXDRVTRIM_HS_0DB_M2(6'b011011), .PMA_SER_DRV_CTRL_M3_TXDRVTRIM_FS_3P5DB_M3(6'b010100)
        , .PMA_SER_DRV_CTRL_M3_TXDRVTRIM_FS_6P0DB_M3(6'b011011), .PMA_SER_DRV_CTRL_M3_TXDRVTRIM_HS_0DB_M3(6'b011011)
        , .PMA_SER_DRV_CTRL_M4_TXDRVTRIM_FS_3P5DB_M4(6'b001010), .PMA_SER_DRV_CTRL_M4_TXDRVTRIM_FS_6P0DB_M4(6'b001100)
        , .PMA_SER_DRV_CTRL_M4_TXDRVTRIM_HS_0DB_M4(6'b100100), .PMA_SER_DRV_CTRL_M5_TXDRVTRIM_BEACON_3P5DB_0(6'b111000)
        , .PMA_SER_DRV_CTRL_M5_TXDRVTRIM_BEACON_3P5DB_1(6'b111011), .PMA_SER_DRV_CTRL_M5_TXDRVTRIM_BEACON_6P0DB_0(6'b111000)
        , .PMA_SER_DRV_CTRL_M5_TXDRVTRIM_BEACON_6P0DB_1(6'b011011), .PMA_SERDES_RTL_CTRL_RESET_RTL(1'b0)
        , .PMA_SERDES_RTL_CTRL_TX_PRBSMODE(3'b000), .PMA_SERDES_RTL_CTRL_TX_DATA_SELECT(3'b000)
        , .PMA_SERDES_RTL_CTRL_RX_DATA_SELECT(2'b00), .PMA_SERDES_RTL_CTRL_RX_FIFO_INPUT_SELECT_NEIGHBOR(1'b0)
        , .PMA_SERDES_RTL_CTRL_RX_EYEMONITOR_COMPARISON_DATA_SEL(1'b0)
        , .PMA_DES_DFE_CAL_CTRL_0_DFE_CAL_CEN(1'b0), .PMA_DES_DFE_CAL_CTRL_0_DFE_CAL_RESET(1'b1)
        , .PMA_DES_DFE_CAL_CTRL_0_EN_FE_CAL(1'b0), .PMA_DES_DFE_CAL_CTRL_0_EN_DFE_CAL(1'b0)
        , .PMA_DES_DFE_CAL_CTRL_0_EN_OFFSET_CAL(1'b0), .PMA_DES_DFE_CAL_CTRL_0_WAIT_PERIOD_GOOD_LOCK(3'b111)
        , .PMA_DES_DFE_CAL_CTRL_0_NUM_SAMPLES_CTLE_OFFSET_CAL(6'b010000)
        , .PMA_DES_DFE_CAL_CTRL_0_NUM_SAMPLES_GOOD_LOCK(8'b01100100), .PMA_DES_DFE_CAL_CTRL_1_BYPASS_DFECAL_USER(1'b0)
        , .PMA_DES_DFE_CAL_CTRL_1_DFE_CAL_EM_ONLY(1'b0), .PMA_DES_DFE_CAL_CTRL_1_DFE_CAL_FORCEH(1'b0)
        , .PMA_DES_DFE_CAL_CTRL_1_PHASE_DIRECTION_USER(1'b1), .PMA_DES_DFE_CAL_CTRL_1_DFE_CAL_CLKDIV(4'b0001)
        , .PMA_DES_DFE_CAL_CTRL_1_DFE_CAL_FREQUENCY(3'b000), .PMA_DES_DFE_CAL_CTRL_1_DFE_CAL_FORCE_CDR_COEFFS(1'b0)
        , .PMA_DES_DFE_CAL_CTRL_1_DFE_CAL_NUM_COEFFS(3'b100), .PMA_DES_DFE_CAL_CTRL_1_MAX_DFE_CYCLES(5'b00011)
        , .PMA_DES_DFE_CAL_CTRL_1_MAX_AREA_CYCLES(2'b01), .PMA_DES_DFE_CAL_CTRL_2_SETALT_OFFSET_DFE0(1'b0)
        , .PMA_DES_DFE_CAL_CTRL_2_SETALT_OFFSET_DFE1(1'b0), .PMA_DES_DFE_CAL_CTRL_2_SETALT_OFFSET_EM0(1'b0)
        , .PMA_DES_DFE_CAL_CTRL_2_SETALT_OFFSET_EM1(1'b0), .PMA_DES_DFE_CAL_CTRL_2_SET_DFE_COEFFS_USER(1'b0)
        , .PMA_DES_DFE_CAL_CTRL_2_ERROR_THR_CHANNEL_ALIGN(12'b000010000000)
        , .PMA_DES_DFE_CAL_CMD_RUN_CTLE_OFFSET_CAL0_USER(1'b0), .PMA_DES_DFE_CAL_CMD_RUN_CTLE_OFFSET_CAL1_USER(1'b0)
        , .PMA_DES_DFE_CAL_CMD_RUN_CTLE_OFFSET_CAL2_USER(1'b0), .PMA_DES_DFE_CAL_CMD_RUN_CTLE_OFFSET_CAL3_USER(1'b0)
        , .PMA_DES_DFE_CAL_CMD_RUN_CTLE_OFFSET_CAL4_USER(1'b0), .PMA_DES_DFE_CAL_CMD_RUN_CTLE_OFFSET_CAL5_USER(1'b0)
        , .PMA_DES_DFE_CAL_CMD_RUN_CTLE_OFFSET_CAL6_USER(1'b0), .PMA_DES_DFE_CAL_CMD_RUN_CTLE_OFFSET_CAL7_USER(1'b0)
        , .PMA_DES_DFE_CAL_CMD_RUN_AREA_COMPUTE_USER(1'b0), .PMA_DES_DFE_CAL_CMD_RUN_CHANNEL_ALIGN_USER(1'b0)
        , .PMA_DES_DFE_CAL_CMD_RUN_CENTER_HORIZONTAL_EM_USER(1'b0), .PMA_DES_DFE_CAL_CMD_RUN_CENTER_HORIZONTAL_USER(1'b0)
        , .PMA_DES_DFE_CAL_CMD_RUN_HORIZONTAL_EM_USER(1'b0), .PMA_DES_DFE_CAL_CMD_RUN_HORIZONTAL_USER(1'b0)
        , .PMA_DES_DFE_CAL_CMD_RUN_VERTICAL_EM_USER(1'b0), .PMA_DES_DFE_CAL_CMD_RUN_VERTICAL_USER(1'b0)
        , .PMA_DES_DFE_CAL_CMD_RUN_DFECAL_USER(1'b0), .PMA_DES_DFE_CAL_CMD_RUN_FE_CALIBRATION_USER(1'b0)
        , .PMA_DES_DFE_CAL_CMD_RUN_FULL_CAL_USER(1'b0), .PMA_DES_DFE_CAL_CMD_RUN_GOOD_LOCK_USER(1'b0)
        , .PMA_DES_DFE_CAL_CMD_RUN_STEP_PHASE_DFE_USER(1'b0), .PMA_DES_DFE_CAL_CMD_RUN_STEP_PHASE_EM_USER(1'b0)
        , .PMA_DES_DFE_CAL_BYPASS_SEL_H0CDR(1'b0), .PMA_DES_DFE_CAL_BYPASS_SEL_H0DFE(1'b0)
        , .PMA_DES_DFE_CAL_BYPASS_SEL_H0EM(1'b0), .PMA_DES_DFE_CAL_BYPASS_SEL_H1(1'b0)
        , .PMA_DES_DFE_CAL_BYPASS_SEL_H2(1'b0), .PMA_DES_DFE_CAL_BYPASS_SEL_H3(1'b0)
        , .PMA_DES_DFE_CAL_BYPASS_SEL_H4(1'b0), .PMA_DES_DFE_CAL_BYPASS_SEL_H5(1'b0)
        , .PMA_DES_DFE_CAL_BYPASS_SEL_CALIBRATION_CLK_EN(1'b0), .PMA_DES_DFE_CAL_BYPASS_SEL_CDRCTLE(1'b0)
        , .PMA_DES_DFE_CAL_BYPASS_SEL_CST1_DFEEM(1'b0), .PMA_DES_DFE_CAL_BYPASS_SEL_CST2_DFEEM(1'b0)
        , .PMA_DES_DFE_CAL_BYPASS_SEL_CTLEEN_DFE(1'b0), .PMA_DES_DFE_CAL_BYPASS_SEL_CTLEEN_EM(1'b0)
        , .PMA_DES_DFE_CAL_BYPASS_SEL_PHICTRL_DFE(1'b0), .PMA_DES_DFE_CAL_BYPASS_SEL_PHICTRL_EM(1'b0)
        , .PMA_DES_DFE_CAL_BYPASS_SEL_RCVEN(1'b0), .PMA_DES_DFE_CAL_BYPASS_SEL_RST1_DFEEM(1'b0)
        , .PMA_DES_DFE_CAL_BYPASS_SEL_RST2_DFEEM(1'b0), .PMA_DES_DFE_CAL_BYPASS_SEL_RUN_EYEMONITOR_COMPARISON(1'b0)
        , .PMA_DES_DFE_CAL_BYPASS_SEL_SLIP_DES_EM(1'b0), .PMA_DES_DFE_CAL_BYPASS_SEL_LOCK_OVERRIDE(1'b0)
        , .PCSCMN_SOFT_RESET_NV_MAP(1'b0), .PCSCMN_SOFT_RESET_V_MAP(1'b0)
        , .PCSCMN_SOFT_RESET_PERIPH(1'b0), .PCSCMN_GSSCLK_CTRL_MCLK_GSSCLK_0_SEL(5'b00000)
        , .PCSCMN_GSSCLK_CTRL_MCLK_GSSCLK_1_SEL(5'b00000), .PCSCMN_GSSCLK_CTRL_MCLK_GSSCLK_2_SEL(5'b00000)
        , .PCSCMN_QRST_R0_QRST0_LANE(2'b00), .PCSCMN_QRST_R0_QRST0_RST_SEL(4'b0000)
        , .PCSCMN_QRST_R0_QRST1_LANE(2'b00), .PCSCMN_QRST_R0_QRST1_RST_SEL(4'b0000)
        , .PCSCMN_QDBG_R0_PCS_DBG_MODE(3'b000), .PCSCMN_QDBG_R0_PCS_DBG_LANE_X(2'b00)
        , .PCSCMN_QDBG_R0_PCS_DBG_LANE_Y(2'b01), .PCS_SOFT_RESET_NV_MAP(1'b0)
        , .PCS_SOFT_RESET_V_MAP(1'b0), .PCS_LFWF_R0_RXFWF_WMARK(1'b0)
        , .PCS_LFWF_R0_TXFWF_WMARK(1'b0), .PCS_LPIP_R0_PIPE_SHAREDPLL(1'b1)
        , .PCS_LPIP_R0_PIPE_INITIALIZATION_DONE(1'b1), .PCS_LPIP_R0_PIPE_OOB_IDLEBURST_TIMING(2'b10)
        , .PCS_L64_R0_L64_CFG_BER_1US_TIMER_VAL(11'b00000000000), .PCS_L64_R1_L64_BYPASS_TEST(1'b1)
        , .PCS_L64_R1_L64_CFG_TEST_PATTERN_EN(1'b0), .PCS_L64_R1_L64_CFG_TEST_PATT_TYPE_SEL(1'b0)
        , .PCS_L64_R1_L64_CFG_TEST_PRBS31_EN(1'b0), .PCS_L64_R1_L64_CFG_TEST_PATT_DATA_SEL(1'b0)
        , .PCS_L64_R2_L64_SEED_A_VALUE_LO32(32'b00000000000000000000000000000000)
        , .PCS_L64_R3_L64_SEED_A_VALUE_HI26(26'b00000000000000000000000000)
        , .PCS_L64_R4_L64_SEED_B_VALUE_LO32(32'b00000000000000000000000000000000)
        , .PCS_L64_R5_L64_SEED_B_VALUE_HI26(26'b00000000000000000000000000)
        , .PCS_L64_R6_L64_TX_ADV_CYC_DLY(5'b00000), .PCS_L64_R6_L64_TX_ADD_UI(16'b0000000000000000)
        , .PCS_L64_R7_L64_RX_ADV_CYC_DLY(5'b00000), .PCS_L64_R7_L64_RX_ADD_UI(16'b0000000000000000)
        , .PCS_L8_R0_L8_TXENCSWAPSEL(1'b0), .PCS_LRST_R0_LRST_SOFT_PCS_RX_RESET(1'b0)
        , .PCS_LRST_R0_LRST_SOFT_PCS_RX_DIV2_RESET(1'b0), .PCS_LRST_R0_LRST_ULCKD_CDR_RESETS_PCS_RX(1'b1)
        , .PCS_LRST_R0_LRST_SOFT_RXFWF_RESET(1'b0), .PCS_LRST_R0_LRST_SOFT_PCS_TX_RESET(1'b0)
        , .PCS_LRST_R0_LRST_SOFT_PCS_TX_DIV2_RESET(1'b0), .PCS_LRST_R0_LRST_ULCKD_PLL_RESETS_PCS_TX(1'b0)
        , .PCS_LRST_R0_LRST_SOFT_TXFWF_RESET(1'b0), .PCS_LRST_R0_LRST_SOFT_PIPE_RESET(7'b0000000)
        , .PCS_LRST_OPT_LRST_DISABLE_FAB_PCS_RESET_FOR_RX(1'b0), .PCS_LRST_OPT_LRST_DISABLE_FAB_PCS_RESET_FOR_TX(1'b0)
        , .PCS_OOB_R0_OOB_BURST_MIN_CYCLE(8'b00001111), .PCS_OOB_R0_OOB_BURST_MAX_CYCLE(8'b00010001)
        , .PCS_OOB_R0_OOB_WAKE_MIN_CYCLE(8'b00001111), .PCS_OOB_R0_OOB_WAKE_MAX_CYCLE(8'b00010001)
        , .PCS_OOB_R1_OOB_RST_INIT_MIN_CYCLE(8'b00101101), .PCS_OOB_R1_OOB_RST_INIT_MAX_CYCLE(8'b00110011)
        , .PCS_OOB_R1_OOB_SAS_MIN_CYCLE(8'b10001000), .PCS_OOB_R1_OOB_SAS_MAX_CYCLE(8'b10011000)
        , .PCS_OOB_R2_TXOOB_PROG_DATA_L32B(32'b00000000000000000000000000000000)
        , .PCS_OOB_R3_TXOOB_PROG_DATA_H8B(8'b00000000), .PCS_PMA_CTRL_R0_PMA_P2_ENTER_INT_MASK(1'b1)
        , .PCS_PMA_CTRL_R0_PMA_P2_EXIT_INT_MASK(1'b1), .PCS_PMA_CTRL_R0_PMA_P2_ENTER_INT(1'b0)
        , .PCS_PMA_CTRL_R0_PMA_P2_EXIT_INT(1'b0), .PCS_PMA_CTRL_R0_PMA_RXPLL_LOCK_INT_MASK(1'b1)
        , .PCS_PMA_CTRL_R0_PMA_RXPLL_UNLOCK_INT_MASK(1'b1), .PCS_PMA_CTRL_R0_PMA_RXPLL_LOCK_INT(1'b0)
        , .PCS_PMA_CTRL_R0_PMA_RXPLL_UNLOCK_INT(1'b0), .PCS_PMA_CTRL_R0_PMA_RXPLL_FLOCK_SEL(1'b0)
        , .PCS_PMA_CTRL_R0_PMA_TXPLL_LOCK_INT_MASK(1'b1), .PCS_PMA_CTRL_R0_PMA_TXPLL_UNLOCK_INT_MASK(1'b1)
        , .PCS_PMA_CTRL_R0_PMA_TXPLL_LOCK_INT(1'b0), .PCS_PMA_CTRL_R0_PMA_TXPLL_UNLOCK_INT(1'b0)
        , .PCS_PMA_CTRL_R1_RXBEACON_MAX_PULSE_WIDTH(11'b11001000000), .PCS_PMA_CTRL_R1_TXBEACON_PULSE_WIDTH(12'b000000001010)
        , .PCS_PMA_CTRL_R2_PD_PLL_CNT(8'b10100110), .PCS_PMA_CTRL_R2_PIPE_RATE_INIT(2'b00)
        , .PCS_PMA_CTRL_R2_FAB_DRIVES_TXPADS(1'b0), .PCS_MSTR_CTRL_LANE_MSTR(2'b00)
        , .MAIN_SOFT_RESET_PERIPH(1'b0), .MAIN_SOFT_RESET_NV_MAP(1'b0)
        , .MAIN_SOFT_RESET_V_MAP(1'b0), .MAIN_MAJOR_PCIE_USAGE_MODE(4'b1000)
        , .MAIN_INT_PIPE_CLK_CTRL_PCLK_INT_LN0_SEL(2'b10), .MAIN_INT_PIPE_CLK_CTRL_PCLK_INT_LN1_SEL(2'b10)
        , .MAIN_INT_PIPE_CLK_CTRL_PCLK_INT_LN2_SEL(1'b0), .MAIN_INT_PIPE_CLK_CTRL_PCLK_INT_LN3_SEL(1'b1)
        , .MAIN_EXT_PIPE_CLK_CTRL_PCLK_EXT_LN0_SEL(1'b0), .MAIN_EXT_PIPE_CLK_CTRL_PCLK_EXT_LN1_SEL(1'b0)
        , .MAIN_EXT_PIPE_CLK_CTRL_PCLK_EXT_LN2_SEL(1'b0), .MAIN_EXT_PIPE_CLK_CTRL_PCLK_EXT_LN3_SEL(1'b0)
        , .MAIN_QMUX_R0_PCIE_DBG_SEL(3'b111), .MAIN_DLL_CTRL0_PHASE_P(2'b11)
        , .MAIN_DLL_CTRL0_PHASE_S(2'b11), .MAIN_DLL_CTRL0_SEL_P(2'b00)
        , .MAIN_DLL_CTRL0_SEL_S(2'b00), .MAIN_DLL_CTRL0_REF_SEL(1'b0)
        , .MAIN_DLL_CTRL0_FB_SEL(1'b0), .MAIN_DLL_CTRL0_DIV_SEL(1'b0)
        , .MAIN_DLL_CTRL0_ALU_UPD(2'b00), .MAIN_DLL_CTRL0_LOCK_FRC(1'b0)
        , .MAIN_DLL_CTRL0_LOCK_FLT(2'b00), .MAIN_DLL_CTRL0_LOCK_HIGH(4'b1000)
        , .MAIN_DLL_CTRL0_LOCK_LOW(4'b1000), .MAIN_DLL_CTRL1_SET_ALU(8'b00000000)
        , .MAIN_DLL_CTRL1_ADJ_DEL4(7'b0000000), .MAIN_DLL_CTRL1_TEST_S(1'b0)
        , .MAIN_DLL_CTRL1_TEST_RING(1'b0), .MAIN_DLL_CTRL1_INIT_CODE(6'b000000)
        , .MAIN_DLL_CTRL1_RELOCK_FAST(1'b0), .MAIN_DLL_STAT0_RESET(1'b0)
        , .MAIN_DLL_STAT0_PHASE_MOVE_CLK(1'b0), .MAIN_OVRLY_AXI0_IFC_MODE(2'b01)
        , .MAIN_OVRLY_AXI1_IFC_MODE(2'b01), .MAIN_INT_PIPE_CLK_CTRL_PCIE_0_PCLK_SEL(3'b110)
        , .MAIN_INT_PIPE_CLK_CTRL_PCIE_1_PCLK_SEL(3'b010), .MAIN_CLK_CTRL_AXI0_CLKENA(1'b0)
        , .MAIN_CLK_CTRL_AXI1_CLKENA(1'b0), .MAIN_DLL_STAT0_LOCK_INT_EN(1'b0)
        , .MAIN_DLL_STAT0_UNLOCK_INT_EN(1'b0), .MAIN_DLL_STAT0_LOCK_INT(1'b0)
        , .MAIN_DLL_STAT0_UNLOCK_INT(1'b1), .MAIN_TEST_DLL_RING_OSC_ENABLE(1'b0)
        , .MAIN_TEST_DLL_REF_ENABLE(1'b0), .MAIN_SPARE_SCRATCHPAD(8'b00000000)
        , .MAIN_SPARE_SPARE_CTRL(24'b011000000000000000000000), .PMA_SOFT_RESET_PERIPH(1'b0)
        , .PMA_DES_CDR_CTRL_3_CST1_CDR(2'b00), .PMA_DES_CDR_CTRL_3_CST2_CDR(2'b00)
        , .PMA_DES_CDR_CTRL_3_RST1_CDR(2'b00), .PMA_DES_CDR_CTRL_3_RST2_CDR(2'b00)
        , .PMA_DES_CDR_CTRL_3_RXDRV_CDR(2'b00), .PMA_DES_DFEEM_CTRL_3_CST1_DFEEM(2'b00)
        , .PMA_DES_DFEEM_CTRL_3_CST2_DFEEM(2'b00), .PMA_DES_DFEEM_CTRL_3_RST1_DFEEM(2'b00)
        , .PMA_DES_DFEEM_CTRL_3_RST2_DFEEM(2'b00), .PMA_DES_DFE_CTRL_2_RXDRV_DFE(2'b00)
        , .PMA_DES_DFE_CTRL_2_CTLEEN_DFE(1'b0), .PMA_DES_EM_CTRL_2_RXDRV_EM(2'b00)
        , .PMA_DES_EM_CTRL_2_CTLEEN_EM(1'b0), .PMA_DES_IN_TERM_RXRTRIM(4'b0111)
        , .PMA_DES_IN_TERM_RXTEN(1'b0), .PMA_DES_IN_TERM_RXRTRIM_SEL(2'b01)
        , .PMA_DES_IN_TERM_ACCOUPLE_RXVCM_EN(1'b1), .PMA_DES_PKDET_RXPKDETEN(1'b1)
        , .PMA_DES_PKDET_RXPKDETRANGE(1'b0), .PMA_DES_PKDET_RXPKDET_LOW_THRESHOLD(3'b001)
        , .PMA_DES_PKDET_RXPKDET_HIGH_THRESHOLD(3'b010), .PMA_DES_RTL_LOCK_CTRL_LOCK_MODE(1'b0)
        , .PMA_DES_RTL_LOCK_CTRL_LOCK_OVERRIDE(2'b00), .PMA_DES_RTL_LOCK_CTRL_FDET_SAMPLE_PERIODS(5'b00001)
        , .PMA_DES_RXPLL_DIV_RXPLL_FBDIV(8'b00011001), .PMA_DES_RXPLL_DIV_RXPLL_REFDIV(5'b00010)
        , .PMA_DES_RXPLL_DIV_RXPLL_RANGE(2'b01), .PMA_DES_RXPLL_DIV_CDR_GAIN(1'b0)
        , .PMA_DES_TEST_BUS_RXATESTEN(1'b0), .PMA_DES_CLK_CTRL_RXREFCLK_SEL(3'b100)
        , .PMA_DES_CLK_CTRL_DESMODE(3'b111), .PMA_DES_CLK_CTRL_DATALOCKEN(1'b0)
        , .PMA_DES_CLK_CTRL_DATALOCKDIVEN(1'b0), .PMA_SER_CTRL_TXVBGREF_SEL(1'b0)
        , .PMA_SER_CLK_CTRL_TXPOSTDIVEN(1'b0), .PMA_SER_CLK_CTRL_TXPOSTDIV(2'b00)
        , .PMA_SER_CLK_CTRL_TXBITCLKSEL(1'b0), .PMA_SER_CLK_CTRL_SERMODE(3'b111)
        , .PMA_SER_DRV_BYP_BYPASS_VALUE(8'b00000000), .PMA_SER_DRV_BYP_TX_BYPASS_SELECT_RTL(2'b00)
        , .PMA_SER_DRV_BYP_TX_BYPASS_SELECT(1'b0), .PMA_SER_RXDET_CTRL_RXDETECT_STEP_WAIT_COUNT(5'b10000)
        , .PMA_SER_TERM_CTRL_TXCM_LEVEL(2'b00), .PMA_SER_TERM_CTRL_TXTEN(1'b0)
        , .PMA_SER_TERM_CTRL_TXRTRIM_SEL(2'b01), .PMA_SER_TERM_CTRL_TXRTRIM(4'b0111)
        , .PMA_SER_TEST_BUS_TXATESTEN(1'b0), .PMA_SER_DRV_DATA_CTRL_TXDEL(16'b0000000000000000)
        , .PMA_SER_DRV_DATA_CTRL_TXDATA_INV(8'b00000000), .PMA_SER_DRV_CTRL_TXDRVTRIM(24'b000000000000000000000000)
        , .PMA_SER_DRV_CTRL_TXDRV(3'b001), .PMA_SER_DRV_CTRL_TXITRIM(2'b10)
        , .PMA_SER_DRV_CTRL_TXODRV(2'b00), .PMA_SER_DRV_CTRL_SEL_TXDRV_CTRL_SEL(1'b0)
        , .PMA_SER_DRV_CTRL_SEL_TXODRV_BOOSTER(1'b0), .PMA_SER_DRV_CTRL_SEL_TXMARGIN(3'b000)
        , .PMA_SER_DRV_CTRL_SEL_TXSWING(1'b0), .PMA_SER_DRV_CTRL_SEL_TXDEEMPHASIS(1'b0)
        , .PMA_SER_DRV_CTRL_SEL_TXDEEMPHASIS_BEACON(1'b0), .PMA_SERDES_RTL_CTRL_RX_HALF_RATE10BIT(1'b0)
        , .PMA_SERDES_RTL_CTRL_TX_HALF_RATE10BIT(1'b0), .PCS_SOFT_RESET_PERIPH(1'b0)
        , .PCS_LFWF_R0_RXFWF_RATIO(2'b00), .PCS_LFWF_R0_TXFWF_RATIO(2'b00)
        , .PCS_LOVR_R0_FAB_IFC_MODE(4'b0000), .PCS_LOVR_R0_PCSPMA_IFC_MODE(4'b0001)
        , .PCS_LPIP_R0_PIPEENABLE(1'b1), .PCS_LPIP_R0_PIPEMODE(1'b0), .PCS_LPIP_R0_PIPE_PCIE_HC(1'b1)
        , .PCS_L64_R0_L64_CFG_BYPASS_SCRAMBLER(1'b0), .PCS_L64_R0_L64_CFG_BYPASS_DISPARITY(1'b1)
        , .PCS_L64_R0_L64_CFG_BYPASS_GEARBOX(1'b0), .PCS_L64_R0_L64_CFG_GRBX_64B67B(1'b0)
        , .PCS_L64_R0_L64_CFG_BER_MON_EN(1'b1), .PCS_L64_R0_L64_CFG_BYPASS_8B_MODE(1'b0)
        , .PCS_L64_R0_L64_CFG_GRBX_SM_C49(1'b0), .PCS_L64_R0_L64_CFG_GRBX_SM_C82(1'b0)
        , .PCS_L8_R0_L8_GEARMODE(2'b00), .PCS_LNTV_R0_LNTV_RX_GEAR(1'b0)
        , .PCS_LNTV_R0_LNTV_RX_IN_WIDTH(3'b111), .PCS_LNTV_R0_LNTV_RX_MODE(1'b0)
        , .PCS_LNTV_R0_LNTV_TX_GEAR(1'b0), .PCS_LNTV_R0_LNTV_TX_OUT_WIDTH(3'b111)
        , .PCS_LNTV_R0_LNTV_TX_MODE(1'b0), .PCS_LCLK_R0_LCLK_EPCS_RX_CLK_SEL(2'b00)
        , .PCS_LCLK_R0_LCLK_EPCS_TX_CLK_SEL(2'b00), .PCS_LCLK_R0_LCLK_TXFWF_TMG_MODE(1'b0)
        , .PCS_LCLK_R0_LCLK_PCS_RX_CLK_SEL(2'b11), .PCS_LCLK_R0_LCLK_PCS_TX_CLK_SEL(2'b11)
        , .PCS_LCLK_R0_LCLK_RXFWF_WCLK_SEL(2'b00), .PCS_LCLK_R0_LCLK_TXFWF_RCLK_SEL(2'b00)
        , .PCS_LCLK_R0_LCLK_RXFWF_WCLK_PIPE(1'b0), .PCS_LCLK_R1_LCLK_ENA_64B6XB_RX_CLK(1'b0)
        , .PCS_LCLK_R1_LCLK_ENA_64B6XB_RX_CLK_DIV2(1'b0), .PCS_LCLK_R1_LCLK_ENA_64B6XB_TX_CLK(1'b0)
        , .PCS_LCLK_R1_LCLK_ENA_64B6XB_TX_CLK_DIV2(1'b0), .PCS_LCLK_R1_LCLK_ENA_8B10B_RX_CLK(1'b0)
        , .PCS_LCLK_R1_LCLK_ENA_8B10B_RXFWF_WCLK(1'b0), .PCS_LCLK_R1_LCLK_ENA_8B10B_TX_CLK(1'b0)
        , .PCS_LCLK_R1_LCLK_ENA_8B10B_TXFWF_RCLK(1'b0), .PCS_LCLK_R1_LCLK_ENA_NATIVE_RX_CLK(1'b0)
        , .PCS_LCLK_R1_LCLK_ENA_NATIVE_RXFWF_WCLK(1'b0), .PCS_LCLK_R1_LCLK_ENA_NATIVE_TX_CLK(1'b0)
        , .PCS_LCLK_R1_LCLK_ENA_NATIVE_TXFWF_RCLK(1'b0), .PCS_LCLK_R1_LCLK_ENA_PIPE_LCL(1'b1)
        , .PCS_LCLK_R1_LCLK_ENA_PIPE_OUT(1'b1), .PCS_PMA_CTRL_R0_PIPE_P0S_EN(1'b1)
        , .PCS_PMA_CTRL_R0_PIPE_P1_EN(1'b1), .PCS_PMA_CTRL_R0_PIPE_P2_EN(1'b1)
        , .PCS_PMA_CTRL_R0_FLASH_FREEZE_P0S_EN(1'b0), .PCS_PMA_CTRL_R0_FLASH_FREEZE_P1_EN(1'b0)
        , .PCS_PMA_CTRL_R0_FLASH_FREEZE_P2_EN(1'b0), .PCS_PMA_CTRL_R0_FAB_EPCS_PMA_RESET_B_EN(1'b1)
         )  PCIESS_LANE3_Pipe_AXI0 (.M_AWADDR_31(
        PCIESS_AXI_1_M_AWADDR[31]), .M_AWADDR_30(
        PCIESS_AXI_1_M_AWADDR[30]), .M_AWADDR_29(
        PCIESS_AXI_1_M_AWADDR[29]), .M_AWADDR_28(
        PCIESS_AXI_1_M_AWADDR[28]), .M_AWADDR_0(
        PCIESS_AXI_1_M_AWADDR[0]), .M_AWADDR_1(
        PCIESS_AXI_1_M_AWADDR[1]), .M_AWADDR_2(
        PCIESS_AXI_1_M_AWADDR[2]), .M_AWADDR_3(
        PCIESS_AXI_1_M_AWADDR[3]), .M_AWADDR_4(
        PCIESS_AXI_1_M_AWADDR[4]), .M_AWADDR_5(
        PCIESS_AXI_1_M_AWADDR[5]), .M_AWADDR_6(
        PCIESS_AXI_1_M_AWADDR[6]), .M_AWADDR_7(
        PCIESS_AXI_1_M_AWADDR[7]), .M_AWADDR_8(
        PCIESS_AXI_1_M_AWADDR[8]), .M_AWADDR_9(
        PCIESS_AXI_1_M_AWADDR[9]), .M_AWADDR_10(
        PCIESS_AXI_1_M_AWADDR[10]), .M_AWADDR_11(
        PCIESS_AXI_1_M_AWADDR[11]), .M_AWADDR_12(
        PCIESS_AXI_1_M_AWADDR[12]), .M_AWADDR_13(
        PCIESS_AXI_1_M_AWADDR[13]), .M_AWADDR_14(
        PCIESS_AXI_1_M_AWADDR[14]), .M_AWADDR_15(
        PCIESS_AXI_1_M_AWADDR[15]), .M_AWADDR_16(
        PCIESS_AXI_1_M_AWADDR[16]), .M_AWADDR_17(
        PCIESS_AXI_1_M_AWADDR[17]), .M_AWADDR_18(
        PCIESS_AXI_1_M_AWADDR[18]), .M_AWADDR_19(
        PCIESS_AXI_1_M_AWADDR[19]), .M_AWADDR_20(
        PCIESS_AXI_1_M_AWADDR[20]), .M_AWADDR_21(
        PCIESS_AXI_1_M_AWADDR[21]), .M_AWADDR_22(
        PCIESS_AXI_1_M_AWADDR[22]), .M_AWADDR_23(
        PCIESS_AXI_1_M_AWADDR[23]), .M_WDATA({PCIESS_AXI_1_M_WDATA[63], 
        PCIESS_AXI_1_M_WDATA[62], PCIESS_AXI_1_M_WDATA[61], 
        PCIESS_AXI_1_M_WDATA[60], PCIESS_AXI_1_M_WDATA[59], 
        PCIESS_AXI_1_M_WDATA[58], PCIESS_AXI_1_M_WDATA[57], 
        PCIESS_AXI_1_M_WDATA[56], PCIESS_AXI_1_M_WDATA[55], 
        PCIESS_AXI_1_M_WDATA[54], PCIESS_AXI_1_M_WDATA[53], 
        PCIESS_AXI_1_M_WDATA[52], PCIESS_AXI_1_M_WDATA[51], 
        PCIESS_AXI_1_M_WDATA[50], PCIESS_AXI_1_M_WDATA[49], 
        PCIESS_AXI_1_M_WDATA[48], PCIESS_AXI_1_M_WDATA[47], 
        PCIESS_AXI_1_M_WDATA[46], PCIESS_AXI_1_M_WDATA[45], 
        PCIESS_AXI_1_M_WDATA[44], PCIESS_AXI_1_M_WDATA[43], 
        PCIESS_AXI_1_M_WDATA[42], PCIESS_AXI_1_M_WDATA[41], 
        PCIESS_AXI_1_M_WDATA[40], PCIESS_AXI_1_M_WDATA[39], 
        PCIESS_AXI_1_M_WDATA[38], PCIESS_AXI_1_M_WDATA[37], 
        PCIESS_AXI_1_M_WDATA[36], PCIESS_AXI_1_M_WDATA[35], 
        PCIESS_AXI_1_M_WDATA[34], PCIESS_AXI_1_M_WDATA[33], 
        PCIESS_AXI_1_M_WDATA[32], PCIESS_AXI_1_M_WDATA[31], 
        PCIESS_AXI_1_M_WDATA[30], PCIESS_AXI_1_M_WDATA[29], 
        PCIESS_AXI_1_M_WDATA[28], PCIESS_AXI_1_M_WDATA[27], 
        PCIESS_AXI_1_M_WDATA[26], PCIESS_AXI_1_M_WDATA[25], 
        PCIESS_AXI_1_M_WDATA[24], PCIESS_AXI_1_M_WDATA[23], 
        PCIESS_AXI_1_M_WDATA[22], PCIESS_AXI_1_M_WDATA[21], 
        PCIESS_AXI_1_M_WDATA[20], PCIESS_AXI_1_M_WDATA[19], 
        PCIESS_AXI_1_M_WDATA[18], PCIESS_AXI_1_M_WDATA[17], 
        PCIESS_AXI_1_M_WDATA[16], PCIESS_AXI_1_M_WDATA[15], 
        PCIESS_AXI_1_M_WDATA[14], PCIESS_AXI_1_M_WDATA[13], 
        PCIESS_AXI_1_M_WDATA[12], PCIESS_AXI_1_M_WDATA[11], 
        PCIESS_AXI_1_M_WDATA[10], PCIESS_AXI_1_M_WDATA[9], 
        PCIESS_AXI_1_M_WDATA[8], PCIESS_AXI_1_M_WDATA[7], 
        PCIESS_AXI_1_M_WDATA[6], PCIESS_AXI_1_M_WDATA[5], 
        PCIESS_AXI_1_M_WDATA[4], PCIESS_AXI_1_M_WDATA[3], 
        PCIESS_AXI_1_M_WDATA[2], PCIESS_AXI_1_M_WDATA[1], 
        PCIESS_AXI_1_M_WDATA[0]}), .RX_REF_CLK(gnd_net), .M_RDATA({
        PCIESS_AXI_1_M_RDATA[63], PCIESS_AXI_1_M_RDATA[62], 
        PCIESS_AXI_1_M_RDATA[61], PCIESS_AXI_1_M_RDATA[60], 
        PCIESS_AXI_1_M_RDATA[59], PCIESS_AXI_1_M_RDATA[58], 
        PCIESS_AXI_1_M_RDATA[57], PCIESS_AXI_1_M_RDATA[56], 
        PCIESS_AXI_1_M_RDATA[55], PCIESS_AXI_1_M_RDATA[54], 
        PCIESS_AXI_1_M_RDATA[53], PCIESS_AXI_1_M_RDATA[52], 
        PCIESS_AXI_1_M_RDATA[51], PCIESS_AXI_1_M_RDATA[50], 
        PCIESS_AXI_1_M_RDATA[49], PCIESS_AXI_1_M_RDATA[48], 
        PCIESS_AXI_1_M_RDATA[47], PCIESS_AXI_1_M_RDATA[46], 
        PCIESS_AXI_1_M_RDATA[45], PCIESS_AXI_1_M_RDATA[44], 
        PCIESS_AXI_1_M_RDATA[43], PCIESS_AXI_1_M_RDATA[42], 
        PCIESS_AXI_1_M_RDATA[41], PCIESS_AXI_1_M_RDATA[40], 
        PCIESS_AXI_1_M_RDATA[39], PCIESS_AXI_1_M_RDATA[38], 
        PCIESS_AXI_1_M_RDATA[37], PCIESS_AXI_1_M_RDATA[36], 
        PCIESS_AXI_1_M_RDATA[35], PCIESS_AXI_1_M_RDATA[34], 
        PCIESS_AXI_1_M_RDATA[33], PCIESS_AXI_1_M_RDATA[32], 
        PCIESS_AXI_1_M_RDATA[31], PCIESS_AXI_1_M_RDATA[30], 
        PCIESS_AXI_1_M_RDATA[29], PCIESS_AXI_1_M_RDATA[28], 
        PCIESS_AXI_1_M_RDATA[27], PCIESS_AXI_1_M_RDATA[26], 
        PCIESS_AXI_1_M_RDATA[25], PCIESS_AXI_1_M_RDATA[24], 
        PCIESS_AXI_1_M_RDATA[23], PCIESS_AXI_1_M_RDATA[22], 
        PCIESS_AXI_1_M_RDATA[21], PCIESS_AXI_1_M_RDATA[20], 
        PCIESS_AXI_1_M_RDATA[19], PCIESS_AXI_1_M_RDATA[18], 
        PCIESS_AXI_1_M_RDATA[17], PCIESS_AXI_1_M_RDATA[16], 
        PCIESS_AXI_1_M_RDATA[15], PCIESS_AXI_1_M_RDATA[14], 
        PCIESS_AXI_1_M_RDATA[13], PCIESS_AXI_1_M_RDATA[12], 
        PCIESS_AXI_1_M_RDATA[11], PCIESS_AXI_1_M_RDATA[10], 
        PCIESS_AXI_1_M_RDATA[9], PCIESS_AXI_1_M_RDATA[8], 
        PCIESS_AXI_1_M_RDATA[7], PCIESS_AXI_1_M_RDATA[6], 
        PCIESS_AXI_1_M_RDATA[5], PCIESS_AXI_1_M_RDATA[4], 
        PCIESS_AXI_1_M_RDATA[3], PCIESS_AXI_1_M_RDATA[2], 
        PCIESS_AXI_1_M_RDATA[1], PCIESS_AXI_1_M_RDATA[0]}), 
        .S_AWADDR_31(PCIESS_AXI_1_S_AWADDR[31]), .S_AWADDR_30(
        PCIESS_AXI_1_S_AWADDR[30]), .S_AWADDR_28(
        PCIESS_AXI_1_S_AWADDR[28]), .S_AWADDR_0(
        PCIESS_AXI_1_S_AWADDR[0]), .S_AWADDR_1(
        PCIESS_AXI_1_S_AWADDR[1]), .S_AWADDR_2(
        PCIESS_AXI_1_S_AWADDR[2]), .S_AWADDR_3(
        PCIESS_AXI_1_S_AWADDR[3]), .S_AWADDR_4(
        PCIESS_AXI_1_S_AWADDR[4]), .S_AWADDR_5(
        PCIESS_AXI_1_S_AWADDR[5]), .S_AWADDR_6(
        PCIESS_AXI_1_S_AWADDR[6]), .S_AWADDR_7(
        PCIESS_AXI_1_S_AWADDR[7]), .S_AWADDR_8(
        PCIESS_AXI_1_S_AWADDR[8]), .S_AWADDR_9(
        PCIESS_AXI_1_S_AWADDR[9]), .S_AWADDR_10(
        PCIESS_AXI_1_S_AWADDR[10]), .S_AWADDR_11(
        PCIESS_AXI_1_S_AWADDR[11]), .S_AWADDR_12(
        PCIESS_AXI_1_S_AWADDR[12]), .S_AWADDR_13(
        PCIESS_AXI_1_S_AWADDR[13]), .S_AWADDR_14(
        PCIESS_AXI_1_S_AWADDR[14]), .S_AWADDR_15(
        PCIESS_AXI_1_S_AWADDR[15]), .S_AWADDR_16(
        PCIESS_AXI_1_S_AWADDR[16]), .S_AWADDR_17(
        PCIESS_AXI_1_S_AWADDR[17]), .S_AWADDR_18(
        PCIESS_AXI_1_S_AWADDR[18]), .S_AWADDR_19(
        PCIESS_AXI_1_S_AWADDR[19]), .S_AWADDR_20(
        PCIESS_AXI_1_S_AWADDR[20]), .S_AWADDR_21(
        PCIESS_AXI_1_S_AWADDR[21]), .S_AWADDR_22(
        PCIESS_AXI_1_S_AWADDR[22]), .S_AWADDR_23(
        PCIESS_AXI_1_S_AWADDR[23]), .M_AWADDR_HW_0(
        PCIE_1_M_AWADDR_0_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_0_net), 
        .M_AWADDR_HW_1(
        PCIE_1_M_AWADDR_1_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_1_net), 
        .M_AWADDR_HW_2(
        PCIE_1_M_AWADDR_2_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_2_net), 
        .M_AWADDR_HW_3(
        PCIE_1_M_AWADDR_3_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_3_net), 
        .M_AWADDR_HW_4(
        PCIE_1_M_AWADDR_4_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_4_net), 
        .M_AWADDR_HW_5(
        PCIE_1_M_AWADDR_5_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_5_net), 
        .M_AWADDR_HW_6(
        PCIE_1_M_AWADDR_6_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_6_net), 
        .M_AWADDR_HW_7(
        PCIE_1_M_AWADDR_7_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_7_net), 
        .M_AWADDR_HW_8(
        PCIE_1_M_AWADDR_8_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_8_net), 
        .M_AWADDR_HW_9(
        PCIE_1_M_AWADDR_9_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_9_net), 
        .M_AWADDR_HW_10(
        PCIE_1_M_AWADDR_10_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_10_net), 
        .M_AWADDR_HW_11(
        PCIE_1_M_AWADDR_11_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_11_net), 
        .M_AWADDR_HW_12(
        PCIE_1_M_AWADDR_12_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_12_net), 
        .M_AWADDR_HW_13(
        PCIE_1_M_AWADDR_13_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_13_net), 
        .M_AWADDR_HW_14(
        PCIE_1_M_AWADDR_14_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_14_net), 
        .M_AWADDR_HW_15(
        PCIE_1_M_AWADDR_15_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_15_net), 
        .M_AWADDR_HW_16(
        PCIE_1_M_AWADDR_16_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_16_net), 
        .M_AWADDR_HW_17(
        PCIE_1_M_AWADDR_17_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_17_net), 
        .M_AWADDR_HW_18(
        PCIE_1_M_AWADDR_18_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_18_net), 
        .M_AWADDR_HW_19(
        PCIE_1_M_AWADDR_19_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_19_net), 
        .M_AWADDR_HW_20(
        PCIE_1_M_AWADDR_20_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_20_net), 
        .M_AWADDR_HW_21(
        PCIE_1_M_AWADDR_21_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_21_net), 
        .M_AWADDR_HW_22(
        PCIE_1_M_AWADDR_22_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_22_net), 
        .M_AWADDR_HW_23(
        PCIE_1_M_AWADDR_23_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_23_net), 
        .M_AWADDR_HW_28(
        PCIE_1_M_AWADDR_28_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_28_net), 
        .M_AWADDR_HW_29(
        PCIE_1_M_AWADDR_29_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_29_net), 
        .M_AWADDR_HW_30(
        PCIE_1_M_AWADDR_30_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_30_net), 
        .M_AWADDR_HW_31(
        PCIE_1_M_AWADDR_31_PCIESS_LANE3_Pipe_AXI0_M_AWADDR_HW_31_net), 
        .M_RDATA_HW({
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_63, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_62, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_61, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_60, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_59, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_58, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_57, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_56, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_55, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_54, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_53, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_52, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_51, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_50, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_49, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_48, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_47, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_46, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_45, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_44, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_43, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_42, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_41, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_40, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_39, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_38, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_37, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_36, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_35, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_34, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_33, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_32, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_31, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_30, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_29, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_28, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_27, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_26, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_25, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_24, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_23, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_22, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_21, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_20, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_19, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_18, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_17, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_16, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_15, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_14, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_13, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_12, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_11, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_10, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_9, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_8, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_7, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_6, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_5, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_4, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_3, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_2, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_1, 
        PCIE_1_M_RDATA_PCIESS_LANE3_Pipe_AXI0_M_RDATA_HW_net_0}), 
        .M_WDATA_HW({
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_63, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_62, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_61, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_60, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_59, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_58, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_57, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_56, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_55, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_54, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_53, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_52, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_51, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_50, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_49, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_48, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_47, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_46, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_45, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_44, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_43, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_42, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_41, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_40, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_39, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_38, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_37, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_36, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_35, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_34, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_33, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_32, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_31, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_30, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_29, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_28, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_27, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_26, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_25, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_24, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_23, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_22, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_21, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_20, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_19, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_18, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_17, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_16, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_15, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_14, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_13, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_12, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_11, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_10, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_9, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_8, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_7, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_6, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_5, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_4, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_3, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_2, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_1, 
        PCIE_1_M_WDATA_PCIESS_LANE3_Pipe_AXI0_M_WDATA_HW_net_0}), 
        .S_AWADDR_HW_0(
        PCIE_1_S_AWADDR_0_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_0_net), 
        .S_AWADDR_HW_1(
        PCIE_1_S_AWADDR_1_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_1_net), 
        .S_AWADDR_HW_2(
        PCIE_1_S_AWADDR_2_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_2_net), 
        .S_AWADDR_HW_3(
        PCIE_1_S_AWADDR_3_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_3_net), 
        .S_AWADDR_HW_4(
        PCIE_1_S_AWADDR_4_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_4_net), 
        .S_AWADDR_HW_5(
        PCIE_1_S_AWADDR_5_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_5_net), 
        .S_AWADDR_HW_6(
        PCIE_1_S_AWADDR_6_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_6_net), 
        .S_AWADDR_HW_7(
        PCIE_1_S_AWADDR_7_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_7_net), 
        .S_AWADDR_HW_8(
        PCIE_1_S_AWADDR_8_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_8_net), 
        .S_AWADDR_HW_9(
        PCIE_1_S_AWADDR_9_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_9_net), 
        .S_AWADDR_HW_10(
        PCIE_1_S_AWADDR_10_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_10_net), 
        .S_AWADDR_HW_11(
        PCIE_1_S_AWADDR_11_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_11_net), 
        .S_AWADDR_HW_12(
        PCIE_1_S_AWADDR_12_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_12_net), 
        .S_AWADDR_HW_13(
        PCIE_1_S_AWADDR_13_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_13_net), 
        .S_AWADDR_HW_14(
        PCIE_1_S_AWADDR_14_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_14_net), 
        .S_AWADDR_HW_15(
        PCIE_1_S_AWADDR_15_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_15_net), 
        .S_AWADDR_HW_16(
        PCIE_1_S_AWADDR_16_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_16_net), 
        .S_AWADDR_HW_17(
        PCIE_1_S_AWADDR_17_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_17_net), 
        .S_AWADDR_HW_18(
        PCIE_1_S_AWADDR_18_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_18_net), 
        .S_AWADDR_HW_19(
        PCIE_1_S_AWADDR_19_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_19_net), 
        .S_AWADDR_HW_20(
        PCIE_1_S_AWADDR_20_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_20_net), 
        .S_AWADDR_HW_21(
        PCIE_1_S_AWADDR_21_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_21_net), 
        .S_AWADDR_HW_22(
        PCIE_1_S_AWADDR_22_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_22_net), 
        .S_AWADDR_HW_23(
        PCIE_1_S_AWADDR_23_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_23_net), 
        .S_AWADDR_HW_28(
        PCIE_1_S_AWADDR_28_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_28_net), 
        .S_AWADDR_HW_30(
        PCIE_1_S_AWADDR_30_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_30_net), 
        .S_AWADDR_HW_31(
        PCIE_1_S_AWADDR_31_PCIESS_LANE3_Pipe_AXI0_S_AWADDR_HW_31_net), 
        .PCS_DEBUG({
        PCIE_COMMON_INSTANCE_PCS_DEBUG_3_PCIESS_LANE3_Pipe_AXI0_PCS_DEBUG_net_19, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_3_PCIESS_LANE3_Pipe_AXI0_PCS_DEBUG_net_18, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_3_PCIESS_LANE3_Pipe_AXI0_PCS_DEBUG_net_17, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_3_PCIESS_LANE3_Pipe_AXI0_PCS_DEBUG_net_16, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_3_PCIESS_LANE3_Pipe_AXI0_PCS_DEBUG_net_15, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_3_PCIESS_LANE3_Pipe_AXI0_PCS_DEBUG_net_14, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_3_PCIESS_LANE3_Pipe_AXI0_PCS_DEBUG_net_13, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_3_PCIESS_LANE3_Pipe_AXI0_PCS_DEBUG_net_12, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_3_PCIESS_LANE3_Pipe_AXI0_PCS_DEBUG_net_11, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_3_PCIESS_LANE3_Pipe_AXI0_PCS_DEBUG_net_10, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_3_PCIESS_LANE3_Pipe_AXI0_PCS_DEBUG_net_9, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_3_PCIESS_LANE3_Pipe_AXI0_PCS_DEBUG_net_8, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_3_PCIESS_LANE3_Pipe_AXI0_PCS_DEBUG_net_7, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_3_PCIESS_LANE3_Pipe_AXI0_PCS_DEBUG_net_6, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_3_PCIESS_LANE3_Pipe_AXI0_PCS_DEBUG_net_5, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_3_PCIESS_LANE3_Pipe_AXI0_PCS_DEBUG_net_4, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_3_PCIESS_LANE3_Pipe_AXI0_PCS_DEBUG_net_3, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_3_PCIESS_LANE3_Pipe_AXI0_PCS_DEBUG_net_2, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_3_PCIESS_LANE3_Pipe_AXI0_PCS_DEBUG_net_1, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_3_PCIESS_LANE3_Pipe_AXI0_PCS_DEBUG_net_0})
        , .REF_CLK_N(gnd_net), .REF_CLK_P(gnd_net), .RX_N(), .RX_P(), 
        .TX_N(), .TX_P(), .JA_CLK(), .TX_BIT_CLK_0(gnd_net), 
        .TX_BIT_CLK_1(gnd_net), .TX_PLL_LOCK_0(gnd_net), 
        .TX_PLL_LOCK_1(gnd_net), .TX_PLL_REF_CLK_0(gnd_net), 
        .TX_PLL_REF_CLK_1(gnd_net), .TX_CLK_G(), .RX_CLK_G(), 
        .PMA_DEBUG(
        PCIE_COMMON_INSTANCE_PMA_DEBUG_3_PCIESS_LANE3_Pipe_AXI0_PMA_DEBUG_net)
        , .ARST_N({nc306, nc307}), .DRI_CLK(gnd_net), .DRI_CTRL({
        gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, 
        gnd_net, gnd_net, gnd_net, gnd_net}), .DRI_WDATA({gnd_net, 
        gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, 
        gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, 
        gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, 
        gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, 
        gnd_net, gnd_net, gnd_net, gnd_net}), .DRI_ARST_N(vcc_net), 
        .DRI_RDATA({nc308, nc309, nc310, nc311, nc312, nc313, nc314, 
        nc315, nc316, nc317, nc318, nc319, nc320, nc321, nc322, nc323, 
        nc324, nc325, nc326, nc327, nc328, nc329, nc330, nc331, nc332, 
        nc333, nc334, nc335, nc336, nc337, nc338, nc339, nc340}), 
        .DRI_INTERRUPT(), .PHYSTATUS_0(
        PCIE_1_PHYSTATUS_3_PCIESS_LANE3_Pipe_AXI0_PHYSTATUS_0_net), 
        .POWERDOWN({
        PCIE_1_POWERDOWN_PCIESS_LANE2_Pipe_AXI1_POWERDOWN_net_1, 
        PCIE_1_POWERDOWN_PCIESS_LANE2_Pipe_AXI1_POWERDOWN_net_0}), 
        .RATE({PCIE_1_RATE_PCIESS_LANE2_Pipe_AXI1_RATE_net_1, 
        PCIE_1_RATE_PCIESS_LANE2_Pipe_AXI1_RATE_net_0}), .RESET_N(
        PCIE_1_RESET_N_PCIESS_LANE2_Pipe_AXI1_RESET_N_net), .RXDATA_0({
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_31, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_30, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_29, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_28, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_27, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_26, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_25, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_24, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_23, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_22, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_21, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_20, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_19, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_18, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_17, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_16, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_15, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_14, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_13, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_12, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_11, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_10, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_9, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_8, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_7, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_6, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_5, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_4, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_3, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_2, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_1, 
        PCIE_1_RXDATA_3_PCIESS_LANE3_Pipe_AXI0_RXDATA_0_net_0}), 
        .RXDATAK_0({
        PCIE_1_RXDATAK_3_PCIESS_LANE3_Pipe_AXI0_RXDATAK_0_net_3, 
        PCIE_1_RXDATAK_3_PCIESS_LANE3_Pipe_AXI0_RXDATAK_0_net_2, 
        PCIE_1_RXDATAK_3_PCIESS_LANE3_Pipe_AXI0_RXDATAK_0_net_1, 
        PCIE_1_RXDATAK_3_PCIESS_LANE3_Pipe_AXI0_RXDATAK_0_net_0}), 
        .RXELECIDLE_0(
        PCIE_1_RXELECIDLE_3_PCIESS_LANE3_Pipe_AXI0_RXELECIDLE_0_net), 
        .RXPOLARITY_0(
        PCIE_1_RXPOLARITY_3_PCIESS_LANE3_Pipe_AXI0_RXPOLARITY_0_net), 
        .RXSTANDBYSTATUS_0(
        PCIE_1_RXSTANDBYSTATUS_3_PCIESS_LANE3_Pipe_AXI0_RXSTANDBYSTATUS_0_net)
        , .RXSTATUS_0({
        PCIE_1_RXSTATUS_3_PCIESS_LANE3_Pipe_AXI0_RXSTATUS_0_net_2, 
        PCIE_1_RXSTATUS_3_PCIESS_LANE3_Pipe_AXI0_RXSTATUS_0_net_1, 
        PCIE_1_RXSTATUS_3_PCIESS_LANE3_Pipe_AXI0_RXSTATUS_0_net_0}), 
        .RXVALID_0(
        PCIE_1_RXVALID_3_PCIESS_LANE3_Pipe_AXI0_RXVALID_0_net), 
        .TXCOMPLIANCE_0(
        PCIE_1_TXCOMPLIANCE_3_PCIESS_LANE3_Pipe_AXI0_TXCOMPLIANCE_0_net)
        , .TXDATA_0({
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_31, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_30, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_29, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_28, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_27, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_26, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_25, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_24, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_23, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_22, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_21, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_20, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_19, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_18, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_17, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_16, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_15, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_14, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_13, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_12, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_11, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_10, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_9, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_8, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_7, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_6, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_5, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_4, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_3, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_2, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_1, 
        PCIE_1_TXDATA_3_PCIESS_LANE3_Pipe_AXI0_TXDATA_0_net_0}), 
        .TXDATAK_0({
        PCIE_1_TXDATAK_3_PCIESS_LANE3_Pipe_AXI0_TXDATAK_0_net_3, 
        PCIE_1_TXDATAK_3_PCIESS_LANE3_Pipe_AXI0_TXDATAK_0_net_2, 
        PCIE_1_TXDATAK_3_PCIESS_LANE3_Pipe_AXI0_TXDATAK_0_net_1, 
        PCIE_1_TXDATAK_3_PCIESS_LANE3_Pipe_AXI0_TXDATAK_0_net_0}), 
        .TXDATAVALID_0(
        PCIE_1_TXDATAVALID_3_PCIESS_LANE3_Pipe_AXI0_TXDATAVALID_0_net), 
        .TXDEEMPH(PCIE_1_TXDEEMPH_PCIESS_LANE2_Pipe_AXI1_TXDEEMPH_net), 
        .TXDETECTRX_LOOPBACK_0(
        PCIE_1_TXDETECTRX_LOOPBACK_3_PCIESS_LANE3_Pipe_AXI0_TXDETECTRX_LOOPBACK_0_net)
        , .TXELECIDLE_0(
        PCIE_1_TXELECIDLE_3_PCIESS_LANE3_Pipe_AXI0_TXELECIDLE_0_net), 
        .TXMARGIN({
        PCIE_1_TXMARGIN_PCIESS_LANE2_Pipe_AXI1_TXMARGIN_net_2, 
        PCIE_1_TXMARGIN_PCIESS_LANE2_Pipe_AXI1_TXMARGIN_net_1, 
        PCIE_1_TXMARGIN_PCIESS_LANE2_Pipe_AXI1_TXMARGIN_net_0}), 
        .TXSWING(PCIE_1_TXSWING_PCIESS_LANE2_Pipe_AXI1_TXSWING_net), 
        .PIPE_CLK_0(
        PCIE_1_PIPE_CLK_3_PCIESS_LANE3_Pipe_AXI0_PIPE_CLK_0_net), 
        .PCLK_OUT_0(
        PCIE_1_PCLK_OUT_3_PCIESS_LANE3_Pipe_AXI0_PCLK_OUT_0_net), 
        .AXI_CLK(PCIE_COMMON_AXI_CLK_OUT_net), .LINK_CLK(gnd_net), 
        .LINK_ADDR({gnd_net, gnd_net, gnd_net}), .LINK_EN(gnd_net), 
        .LINK_ARST_N(gnd_net), .LINK_WDATA({gnd_net, gnd_net, gnd_net, 
        gnd_net}), .LINK_RDATA({nc341, nc342, nc343, nc344}));
    GND PCIESS_AXI_1_M_AWLEN_6_GndInst (.Y(PCIESS_AXI_1_M_AWLEN[6]));
    GND PCIESS_AXI_1_M_AWBURST_1_GndInst (.Y(PCIESS_AXI_1_M_AWBURST[1])
        );
    XCVR_PIPE_AXI1 #( .MAIN_QMUX_R0_QRST0_SRC(3'b001), .MAIN_QMUX_R0_QRST1_SRC(3'b011)
        , .MAIN_QMUX_R0_QRST2_SRC(3'b000), .MAIN_QMUX_R0_QRST3_SRC(3'b000)
        , .DATA_RATE(5000.0), .REG_FILE(""), .PMA_CMN_SOFT_RESET_NV_MAP(1'b0)
        , .PMA_CMN_SOFT_RESET_V_MAP(1'b0), .PMA_CMN_SOFT_RESET_PERIPH(1'b0)
        , .PMA_CMN_TXPLL_CLKBUF_TXPLL_DUALCLK1_MODE(2'b00), .PMA_CMN_TXPLL_CLKBUF_TXPLL_DUALCLK1_ENTERM(2'b00)
        , .PMA_CMN_TXPLL_CLKBUF_TXPLL_DUALCLK0_MODE(2'b10), .PMA_CMN_TXPLL_CLKBUF_TXPLL_DUALCLK0_ENTERM(2'b00)
        , .PMA_CMN_TXPLL_CLKBUF_TXPLL_DUALCLK1_EN_HYST(1'b0), .PMA_CMN_TXPLL_CLKBUF_TXPLL_DUALCLK0_EN_HYST(1'b0)
        , .PMA_CMN_TXPLL_CLKBUF_TXPLL_CLKBUF_EN_RDIFF(1'b0), .PMA_CMN_TXPLL_CLKBUF_TXPLL_CLKBUF_EN_UDRIVE_P(1'b1)
        , .PMA_CMN_TXPLL_CLKBUF_TXPLL_CLKBUF_EN_UDRIVE_N(1'b1), .PMA_CMN_TXPLL_CLKBUF_TXPLL_CLKBUF_EN_PULLUP(1'b0)
        , .PMA_CMN_TXPLL_CLKBUF_TXPLL_CLKBUF_EN_APAD(1'b0), .PMA_CMN_TXPLL_CTRL_TXPLL_BWSEL(1'b1)
        , .PMA_CMN_TXPLL_CTRL_TXPLL_VBGREF_SEL(1'b0), .PMA_CMN_TXPLL_CTRL_TXPLL_FBDIV_SEL(2'b00)
        , .PMA_CMN_TXPLL_CTRL_TXPLL_DSMPD(1'b0), .PMA_CMN_TXPLL_CTRL_TXPLL_PHASESTEPAMOUNT(8'b00000110)
        , .PMA_CMN_TXPLL_CTRL_TXPLL_STEP_PHASE(1'b0), .PMA_CMN_TXPLL_CTRL_TXPLL_PD(1'b0)
        , .PMA_CMN_TXPLL_CTRL_TXPLL_AUXDIVPD(1'b0), .PMA_CMN_TXPLL_CTRL_TXPLL_CLKRESETEN(1'b0)
        , .PMA_CMN_TXPLL_CTRL_TXPLL_CLKRESET(1'b0), .PMA_CMN_TXPLL_CTRL_RESET_RTL_TXPLL(1'b0)
        , .PMA_CMN_TXPLL_CTRL_RESET_RTL(1'b0), .PMA_CMN_TXPLL_CTRL_TXPLL_FOUTAUXDIV2_SEL(1'b0)
        , .PMA_CMN_TXPLL_CLK_SEL_TXPLL_REFCLK_SEL_HM(2'b11), .PMA_CMN_TXPLL_CLK_SEL_TXPLL_REFCLK_SEL_SM(3'b000)
        , .PMA_CMN_TXPLL_CLK_SEL_CASCADE_CLK_SEL_HM(2'b00), .PMA_CMN_TXPLL_CLK_SEL_CASCADE_CLK_SEL_SM(3'b111)
        , .PMA_CMN_TXPLL_CLK_SEL_TXPLL_JA_FREF_SEL(3'b000), .PMA_CMN_TXPLL_CLK_SEL_CDRCLK_LN01_INT_SEL(3'b111)
        , .PMA_CMN_TXPLL_CLK_SEL_CDRCLK_LN23_INT_SEL(3'b111), .PMA_CMN_TXPLL_CLK_SEL_CDRCLK_OUT_UP_SEL(3'b111)
        , .PMA_CMN_TXPLL_CLK_SEL_CDRCLK_OUT_DN_SEL(3'b111), .PMA_CMN_TXPLL_DIV_1_TXPLL_AUXDIV(12'b000000011001)
        , .PMA_CMN_TXPLL_DIV_1_TXPLL_FBDIV(12'b000000011001), .PMA_CMN_TXPLL_DIV_2_TXPLL_FRAC(24'b000000000000000000000001)
        , .PMA_CMN_TXPLL_DIV_2_TXPLL_REFDIV(6'b000001), .PMA_CMN_TXPLL_JA_1_TXPLL_JA_DIVFIN(16'b0000000001100100)
        , .PMA_CMN_TXPLL_JA_1_TXPLL_JA_DIVFFB(16'b0000000001100100), .PMA_CMN_TXPLL_JA_2_TXPLL_JA_SYNCCNTMAX(32'b00000000000000000000000001100100)
        , .PMA_CMN_TXPLL_JA_3_TXPLL_JA_CNTOFFSET(16'b0000000001100100)
        , .PMA_CMN_TXPLL_JA_3_TXPLL_JA_TARGETCNT(32'b00000000000000000000000001100100)
        , .PMA_CMN_TXPLL_JA_4_TXPLL_JA_OTDLY(16'b0000000000000001), .PMA_CMN_TXPLL_JA_4_TXPLL_JA_FMI(8'b00000001)
        , .PMA_CMN_TXPLL_JA_4_TXPLL_JA_FKI(4'b0001), .PMA_CMN_TXPLL_JA_5_TXPLL_JA_PMP1(8'b00000001)
        , .PMA_CMN_TXPLL_JA_5_TXPLL_JA_PMP2(8'b00000001), .PMA_CMN_TXPLL_JA_5_TXPLL_JA_PMI1(8'b00000001)
        , .PMA_CMN_TXPLL_JA_5_TXPLL_JA_PMI2(8'b00000001), .PMA_CMN_TXPLL_JA_6_TXPLL_JA_PKP1(5'b00001)
        , .PMA_CMN_TXPLL_JA_6_TXPLL_JA_PKP2(5'b00001), .PMA_CMN_TXPLL_JA_6_TXPLL_JA_PKI1(5'b00001)
        , .PMA_CMN_TXPLL_JA_6_TXPLL_JA_PKI2(5'b00001), .PMA_CMN_TXPLL_JA_7_TXPLL_JA_DELAYK(24'b000000000000000000000001)
        , .PMA_CMN_TXPLL_JA_7_TXPLL_JA_FDONLY(1'b1), .PMA_CMN_TXPLL_JA_7_TXPLL_JA_ONTARGETOV(1'b1)
        , .PMA_CMN_TXPLL_JA_7_TXPLL_JA_PROGRAM(1'b1), .PMA_CMN_TXPLL_JA_8_TXPLL_JA_FRAC_PRESET(24'b000000000000000000000000)
        , .PMA_CMN_TXPLL_JA_8_TXPLL_JA_PRESET_EN(1'b0), .PMA_CMN_TXPLL_JA_8_TXPLL_JA_HOLD(1'b0)
        , .PMA_CMN_TXPLL_JA_9_TXPLL_JA_INT_PRESET(12'b000000010100), .PMA_CMN_TXPLL_JA_RST_TXPLL_JA_RESET(1'b1)
        , .PMA_CMN_TXPLL_JA_RST_TXPLL_JA_RESET_FFB_OVERRIDE(1'b0), .PMA_CMN_TXPLL_JA_RST_TXPLL_JA_RESET_FFB_EXT(1'b1)
        , .PMA_CMN_TXPLL_JA_RST_TXPLL_JA_RESET_FIN_OVERRIDE(1'b0), .PMA_CMN_TXPLL_JA_RST_TXPLL_JA_RESET_FIN_EXT(1'b1)
        , .PMA_CMN_TXPLL_JA_RST_TXPLL_JA_RESET_CLKS_OVERRIDE(1'b0), .PMA_CMN_TXPLL_JA_RST_TXPLL_JA_RESET_CLKS_EXT(1'b1)
        , .PMA_CMN_SERDES_SSMOD_SSMOD_DOWNSPREAD(1'b0), .PMA_CMN_SERDES_SSMOD_SSMOD_DISABLE_SSCG(1'b1)
        , .PMA_CMN_SERDES_SSMOD_SSMOD_SPREAD(5'b00000), .PMA_CMN_SERDES_SSMOD_SSMOD_DIVVAL(6'b000001)
        , .PMA_CMN_SERDES_SSMOD_SSMOD_EXT_MAXADDR(8'b01111111), .PMA_CMN_SERDES_SSMOD_SSMOD_SEL_EXTWAVE(2'b00)
        , .PMA_CMN_SERDES_SSMOD_RN_SEL(2'b00), .PMA_CMN_SERDES_SSMOD_RN_FILTER(1'b0)
        , .PMA_CMN_SERDES_RTERM_RTERMCAL85(4'b0011), .PMA_CMN_SERDES_RTERM_RTERMCAL100(4'b0111)
        , .PMA_CMN_SERDES_RTERM_RTERMCAL150(4'b1101), .PMA_CMN_SERDES_RTT_RTT_CAL_TERM(4'b0000)
        , .PMA_CMN_SERDES_RTT_RTT_CURRENT_PROG(2'b00), .PMA_SOFT_RESET_NV_MAP(1'b0)
        , .PMA_SOFT_RESET_V_MAP(1'b0), .PMA_DES_CDR_CTRL_1_DCFBEN_CDR(1'b0)
        , .PMA_DES_CDR_CTRL_1_H0CDR0(5'b00000), .PMA_DES_CDR_CTRL_1_H0CDR1(5'b00000)
        , .PMA_DES_CDR_CTRL_1_H0CDR2(8'b00000000), .PMA_DES_CDR_CTRL_1_H0CDR3(5'b00000)
        , .PMA_DES_CDR_CTRL_1_CMRTRIM_CDR(3'b000), .PMA_DES_CDR_CTRL_2_CSENT1_CDR(2'b01)
        , .PMA_DES_CDR_CTRL_2_CSENT2_CDR(2'b01), .PMA_DES_CDR_CTRL_2_CSENT3_CDR(2'b01)
        , .PMA_DES_CDR_CTRL_3_SLIP_DES_CDR(1'b0), .PMA_DES_CDR_CTRL_3_SLIP_DES_CDR_SEL(1'b0)
        , .PMA_DES_CDR_CTRL_3_SLIP_DES_CDR_EN(1'b0), .PMA_DES_DFEEM_CTRL_1_CSENT1_DFEEM(2'b01)
        , .PMA_DES_DFEEM_CTRL_1_CSENT2_DFEEM(2'b01), .PMA_DES_DFEEM_CTRL_1_CSENT3_DFEEM(2'b01)
        , .PMA_DES_DFEEM_CTRL_1_CMRTRIM_DFEEM(3'b000), .PMA_DES_DFEEM_CTRL_2_H1(5'b00000)
        , .PMA_DES_DFEEM_CTRL_2_H2(5'b00000), .PMA_DES_DFEEM_CTRL_2_H3(5'b00000)
        , .PMA_DES_DFEEM_CTRL_2_H4(5'b00000), .PMA_DES_DFEEM_CTRL_3_H5(5'b00000)
        , .PMA_DES_DFE_CTRL_1_DCFBEN_DFE(1'b0), .PMA_DES_DFE_CTRL_1_H0DFE0(5'b00000)
        , .PMA_DES_DFE_CTRL_1_H0DFE1(5'b00000), .PMA_DES_DFE_CTRL_2_PHICTRL_TH_DFE(8'b00000000)
        , .PMA_DES_DFE_CTRL_2_PHICTRL_GRAY_DFE(3'b000), .PMA_DES_DFE_CTRL_2_SLIP_DES_DFE(1'b0)
        , .PMA_DES_DFE_CTRL_2_SLIP_DES_DFE_SEL(1'b0), .PMA_DES_DFE_CTRL_2_SLIP_DES_DFE_EN(1'b0)
        , .PMA_DES_EM_CTRL_1_DCFBEN_EM(1'b0), .PMA_DES_EM_CTRL_1_H0EM0(5'b00000)
        , .PMA_DES_EM_CTRL_1_H0EM1(5'b00000), .PMA_DES_EM_CTRL_1_CALIBRATION_CLK_EN(1'b0)
        , .PMA_DES_EM_CTRL_2_PHICTRL_TH_EM(8'b00000000), .PMA_DES_EM_CTRL_2_PHICTRL_GRAY_EM(3'b000)
        , .PMA_DES_EM_CTRL_2_SLIP_DES_EM(1'b0), .PMA_DES_EM_CTRL_2_SLIP_DES_EM_SEL(1'b0)
        , .PMA_DES_EM_CTRL_2_SLIP_DES_EM_EN(1'b0), .PMA_DES_RTL_EM_RUN_EYEMONITOR_COMPARISON(1'b0)
        , .PMA_DES_RTL_EM_EYEMONITOR_SAMPLE_COUNT(12'b000001100100), .PMA_DES_RTL_LOCK_CTRL_LOCK_OVERRIDE_FROMFAB(1'b0)
        , .PMA_DES_TEST_BUS_RXATESTSEL(3'b000), .PMA_DES_TEST_BUS_RXDTESTEN(1'b0)
        , .PMA_DES_TEST_BUS_RXDTESTSEL(3'b000), .PMA_DES_CLK_CTRL_RXBYPASSEN(1'b0)
        , .PMA_DES_RSTPD_RXPD(1'b0), .PMA_DES_RSTPD_RESETDES(1'b0), .PMA_DES_RSTPD_PDDFE(1'b1)
        , .PMA_DES_RSTPD_PDEM(1'b1), .PMA_DES_RSTPD_RCVEN(1'b1), .PMA_DES_RSTPD_RESET_FIFO(1'b0)
        , .PMA_DES_RTL_ERR_CHK_READ_ERROR(1'b0), .PMA_DES_PCIE1_2_RXPLL_DIV_PCIE1_RXPLL_FBDIV(8'b00011001)
        , .PMA_DES_PCIE1_2_RXPLL_DIV_PCIE1_RXPLL_REFDIV(5'b00010), .PMA_DES_PCIE1_2_RXPLL_DIV_PCIE1_RXPLL_RANGE(2'b01)
        , .PMA_DES_PCIE1_2_RXPLL_DIV_PCIE2_RXPLL_FBDIV(8'b00110010), .PMA_DES_PCIE1_2_RXPLL_DIV_PCIE2_RXPLL_REFDIV(5'b00010)
        , .PMA_DES_PCIE1_2_RXPLL_DIV_PCIE2_RXPLL_RANGE(2'b00), .PMA_DES_SATA1_2_RXPLL_DIV_SATA1_RXPLL_FBDIV(8'b00011000)
        , .PMA_DES_SATA1_2_RXPLL_DIV_SATA1_RXPLL_REFDIV(5'b00100), .PMA_DES_SATA1_2_RXPLL_DIV_SATA1_RXPLL_RANGE(2'b10)
        , .PMA_DES_SATA1_2_RXPLL_DIV_SATA2_RXPLL_FBDIV(8'b00011000), .PMA_DES_SATA1_2_RXPLL_DIV_SATA2_RXPLL_REFDIV(5'b00010)
        , .PMA_DES_SATA1_2_RXPLL_DIV_SATA2_RXPLL_RANGE(2'b01), .PMA_DES_SATA3_RXPLL_DIV_SATA3_RXPLL_FBDIV(8'b00110000)
        , .PMA_DES_SATA3_RXPLL_DIV_SATA3_RXPLL_REFDIV(5'b00010), .PMA_DES_SATA3_RXPLL_DIV_SATA3_RXPLL_RANGE(2'b00)
        , .PMA_SER_CTRL_CMSTEP_VALUE(1'b0), .PMA_SER_CTRL_CMSTEP(1'b0)
        , .PMA_SER_CTRL_NLPBK_EN(1'b0), .PMA_SER_CTRL_HSLPBKEN(1'b0), .PMA_SER_CTRL_HSLPBK_SEL(3'b000)
        , .PMA_SER_RSTPD_RESETSEREN(1'b1), .PMA_SER_RSTPD_RESETSER(1'b0)
        , .PMA_SER_RSTPD_TXPD(1'b0), .PMA_SER_DRV_BYP_BYPASSSER(1'b0)
        , .PMA_SER_RXDET_CTRL_RXDETECT_COUNT_THRESHOLD(14'b00000000000001)
        , .PMA_SER_RXDET_CTRL_RX_DETECT_EN(1'b0), .PMA_SER_RXDET_CTRL_RXDETECT_START(1'b0)
        , .PMA_SER_STATIC_LSB_STATIC_PATTERN_LSB(20'b00000000000000000000)
        , .PMA_SER_STATIC_MSB_STATIC_PATTERN_MSB(20'b00000000000000000000)
        , .PMA_SER_TEST_BUS_TXATESTSEL(3'b000), .PMA_SER_TEST_BUS_DTESTEN_RTL(1'b0)
        , .PMA_SER_TEST_BUS_DTESTSEL_RTL(4'b0000), .PMA_SER_TEST_BUS_JTAG_TO_DTEST_SEL(3'b000)
        , .PMA_SER_TEST_BUS_PRBSERR_TO_DTEST_SEL(2'b00), .PMA_SER_TEST_BUS_RXPKDETOUT_TO_DTEST_SEL(3'b111)
        , .PMA_SER_DRV_CTRL_M0_TXDRVTRIM_FS_3P5DB_M0(6'b100011), .PMA_SER_DRV_CTRL_M0_TXDRVTRIM_FS_6P0DB_M0(6'b110100)
        , .PMA_SER_DRV_CTRL_M0_TXDRVTRIM_HS_0DB_M0(6'b011011), .PMA_SER_DRV_CTRL_M1_TXDRVTRIM_FS_3P5DB_M1(6'b100111)
        , .PMA_SER_DRV_CTRL_M1_TXDRVTRIM_FS_6P0DB_M1(6'b101100), .PMA_SER_DRV_CTRL_M1_TXDRVTRIM_HS_0DB_M1(6'b100011)
        , .PMA_SER_DRV_CTRL_M2_TXDRVTRIM_FS_3P5DB_M2(6'b011011), .PMA_SER_DRV_CTRL_M2_TXDRVTRIM_FS_6P0DB_M2(6'b011011)
        , .PMA_SER_DRV_CTRL_M2_TXDRVTRIM_HS_0DB_M2(6'b011011), .PMA_SER_DRV_CTRL_M3_TXDRVTRIM_FS_3P5DB_M3(6'b010100)
        , .PMA_SER_DRV_CTRL_M3_TXDRVTRIM_FS_6P0DB_M3(6'b011011), .PMA_SER_DRV_CTRL_M3_TXDRVTRIM_HS_0DB_M3(6'b011011)
        , .PMA_SER_DRV_CTRL_M4_TXDRVTRIM_FS_3P5DB_M4(6'b001010), .PMA_SER_DRV_CTRL_M4_TXDRVTRIM_FS_6P0DB_M4(6'b001100)
        , .PMA_SER_DRV_CTRL_M4_TXDRVTRIM_HS_0DB_M4(6'b100100), .PMA_SER_DRV_CTRL_M5_TXDRVTRIM_BEACON_3P5DB_0(6'b111000)
        , .PMA_SER_DRV_CTRL_M5_TXDRVTRIM_BEACON_3P5DB_1(6'b111011), .PMA_SER_DRV_CTRL_M5_TXDRVTRIM_BEACON_6P0DB_0(6'b111000)
        , .PMA_SER_DRV_CTRL_M5_TXDRVTRIM_BEACON_6P0DB_1(6'b011011), .PMA_SERDES_RTL_CTRL_RESET_RTL(1'b0)
        , .PMA_SERDES_RTL_CTRL_TX_PRBSMODE(3'b000), .PMA_SERDES_RTL_CTRL_TX_DATA_SELECT(3'b000)
        , .PMA_SERDES_RTL_CTRL_RX_DATA_SELECT(2'b00), .PMA_SERDES_RTL_CTRL_RX_FIFO_INPUT_SELECT_NEIGHBOR(1'b0)
        , .PMA_SERDES_RTL_CTRL_RX_EYEMONITOR_COMPARISON_DATA_SEL(1'b0)
        , .PMA_DES_DFE_CAL_CTRL_0_DFE_CAL_CEN(1'b0), .PMA_DES_DFE_CAL_CTRL_0_DFE_CAL_RESET(1'b1)
        , .PMA_DES_DFE_CAL_CTRL_0_EN_FE_CAL(1'b0), .PMA_DES_DFE_CAL_CTRL_0_EN_DFE_CAL(1'b0)
        , .PMA_DES_DFE_CAL_CTRL_0_EN_OFFSET_CAL(1'b0), .PMA_DES_DFE_CAL_CTRL_0_WAIT_PERIOD_GOOD_LOCK(3'b111)
        , .PMA_DES_DFE_CAL_CTRL_0_NUM_SAMPLES_CTLE_OFFSET_CAL(6'b010000)
        , .PMA_DES_DFE_CAL_CTRL_0_NUM_SAMPLES_GOOD_LOCK(8'b01100100), .PMA_DES_DFE_CAL_CTRL_1_BYPASS_DFECAL_USER(1'b0)
        , .PMA_DES_DFE_CAL_CTRL_1_DFE_CAL_EM_ONLY(1'b0), .PMA_DES_DFE_CAL_CTRL_1_DFE_CAL_FORCEH(1'b0)
        , .PMA_DES_DFE_CAL_CTRL_1_PHASE_DIRECTION_USER(1'b1), .PMA_DES_DFE_CAL_CTRL_1_DFE_CAL_CLKDIV(4'b0001)
        , .PMA_DES_DFE_CAL_CTRL_1_DFE_CAL_FREQUENCY(3'b000), .PMA_DES_DFE_CAL_CTRL_1_DFE_CAL_FORCE_CDR_COEFFS(1'b0)
        , .PMA_DES_DFE_CAL_CTRL_1_DFE_CAL_NUM_COEFFS(3'b100), .PMA_DES_DFE_CAL_CTRL_1_MAX_DFE_CYCLES(5'b00011)
        , .PMA_DES_DFE_CAL_CTRL_1_MAX_AREA_CYCLES(2'b01), .PMA_DES_DFE_CAL_CTRL_2_SETALT_OFFSET_DFE0(1'b0)
        , .PMA_DES_DFE_CAL_CTRL_2_SETALT_OFFSET_DFE1(1'b0), .PMA_DES_DFE_CAL_CTRL_2_SETALT_OFFSET_EM0(1'b0)
        , .PMA_DES_DFE_CAL_CTRL_2_SETALT_OFFSET_EM1(1'b0), .PMA_DES_DFE_CAL_CTRL_2_SET_DFE_COEFFS_USER(1'b0)
        , .PMA_DES_DFE_CAL_CTRL_2_ERROR_THR_CHANNEL_ALIGN(12'b000010000000)
        , .PMA_DES_DFE_CAL_CMD_RUN_CTLE_OFFSET_CAL0_USER(1'b0), .PMA_DES_DFE_CAL_CMD_RUN_CTLE_OFFSET_CAL1_USER(1'b0)
        , .PMA_DES_DFE_CAL_CMD_RUN_CTLE_OFFSET_CAL2_USER(1'b0), .PMA_DES_DFE_CAL_CMD_RUN_CTLE_OFFSET_CAL3_USER(1'b0)
        , .PMA_DES_DFE_CAL_CMD_RUN_CTLE_OFFSET_CAL4_USER(1'b0), .PMA_DES_DFE_CAL_CMD_RUN_CTLE_OFFSET_CAL5_USER(1'b0)
        , .PMA_DES_DFE_CAL_CMD_RUN_CTLE_OFFSET_CAL6_USER(1'b0), .PMA_DES_DFE_CAL_CMD_RUN_CTLE_OFFSET_CAL7_USER(1'b0)
        , .PMA_DES_DFE_CAL_CMD_RUN_AREA_COMPUTE_USER(1'b0), .PMA_DES_DFE_CAL_CMD_RUN_CHANNEL_ALIGN_USER(1'b0)
        , .PMA_DES_DFE_CAL_CMD_RUN_CENTER_HORIZONTAL_EM_USER(1'b0), .PMA_DES_DFE_CAL_CMD_RUN_CENTER_HORIZONTAL_USER(1'b0)
        , .PMA_DES_DFE_CAL_CMD_RUN_HORIZONTAL_EM_USER(1'b0), .PMA_DES_DFE_CAL_CMD_RUN_HORIZONTAL_USER(1'b0)
        , .PMA_DES_DFE_CAL_CMD_RUN_VERTICAL_EM_USER(1'b0), .PMA_DES_DFE_CAL_CMD_RUN_VERTICAL_USER(1'b0)
        , .PMA_DES_DFE_CAL_CMD_RUN_DFECAL_USER(1'b0), .PMA_DES_DFE_CAL_CMD_RUN_FE_CALIBRATION_USER(1'b0)
        , .PMA_DES_DFE_CAL_CMD_RUN_FULL_CAL_USER(1'b0), .PMA_DES_DFE_CAL_CMD_RUN_GOOD_LOCK_USER(1'b0)
        , .PMA_DES_DFE_CAL_CMD_RUN_STEP_PHASE_DFE_USER(1'b0), .PMA_DES_DFE_CAL_CMD_RUN_STEP_PHASE_EM_USER(1'b0)
        , .PMA_DES_DFE_CAL_BYPASS_SEL_H0CDR(1'b0), .PMA_DES_DFE_CAL_BYPASS_SEL_H0DFE(1'b0)
        , .PMA_DES_DFE_CAL_BYPASS_SEL_H0EM(1'b0), .PMA_DES_DFE_CAL_BYPASS_SEL_H1(1'b0)
        , .PMA_DES_DFE_CAL_BYPASS_SEL_H2(1'b0), .PMA_DES_DFE_CAL_BYPASS_SEL_H3(1'b0)
        , .PMA_DES_DFE_CAL_BYPASS_SEL_H4(1'b0), .PMA_DES_DFE_CAL_BYPASS_SEL_H5(1'b0)
        , .PMA_DES_DFE_CAL_BYPASS_SEL_CALIBRATION_CLK_EN(1'b0), .PMA_DES_DFE_CAL_BYPASS_SEL_CDRCTLE(1'b0)
        , .PMA_DES_DFE_CAL_BYPASS_SEL_CST1_DFEEM(1'b0), .PMA_DES_DFE_CAL_BYPASS_SEL_CST2_DFEEM(1'b0)
        , .PMA_DES_DFE_CAL_BYPASS_SEL_CTLEEN_DFE(1'b0), .PMA_DES_DFE_CAL_BYPASS_SEL_CTLEEN_EM(1'b0)
        , .PMA_DES_DFE_CAL_BYPASS_SEL_PHICTRL_DFE(1'b0), .PMA_DES_DFE_CAL_BYPASS_SEL_PHICTRL_EM(1'b0)
        , .PMA_DES_DFE_CAL_BYPASS_SEL_RCVEN(1'b0), .PMA_DES_DFE_CAL_BYPASS_SEL_RST1_DFEEM(1'b0)
        , .PMA_DES_DFE_CAL_BYPASS_SEL_RST2_DFEEM(1'b0), .PMA_DES_DFE_CAL_BYPASS_SEL_RUN_EYEMONITOR_COMPARISON(1'b0)
        , .PMA_DES_DFE_CAL_BYPASS_SEL_SLIP_DES_EM(1'b0), .PMA_DES_DFE_CAL_BYPASS_SEL_LOCK_OVERRIDE(1'b0)
        , .PCSCMN_SOFT_RESET_NV_MAP(1'b0), .PCSCMN_SOFT_RESET_V_MAP(1'b0)
        , .PCSCMN_SOFT_RESET_PERIPH(1'b0), .PCSCMN_GSSCLK_CTRL_MCLK_GSSCLK_0_SEL(5'b00000)
        , .PCSCMN_GSSCLK_CTRL_MCLK_GSSCLK_1_SEL(5'b00000), .PCSCMN_GSSCLK_CTRL_MCLK_GSSCLK_2_SEL(5'b00000)
        , .PCSCMN_QRST_R0_QRST0_LANE(2'b00), .PCSCMN_QRST_R0_QRST0_RST_SEL(4'b0000)
        , .PCSCMN_QRST_R0_QRST1_LANE(2'b00), .PCSCMN_QRST_R0_QRST1_RST_SEL(4'b0000)
        , .PCSCMN_QDBG_R0_PCS_DBG_MODE(3'b000), .PCSCMN_QDBG_R0_PCS_DBG_LANE_X(2'b00)
        , .PCSCMN_QDBG_R0_PCS_DBG_LANE_Y(2'b01), .PCS_SOFT_RESET_NV_MAP(1'b0)
        , .PCS_SOFT_RESET_V_MAP(1'b0), .PCS_LFWF_R0_RXFWF_WMARK(1'b0)
        , .PCS_LFWF_R0_TXFWF_WMARK(1'b0), .PCS_LPIP_R0_PIPE_SHAREDPLL(1'b1)
        , .PCS_LPIP_R0_PIPE_INITIALIZATION_DONE(1'b1), .PCS_LPIP_R0_PIPE_OOB_IDLEBURST_TIMING(2'b10)
        , .PCS_L64_R0_L64_CFG_BER_1US_TIMER_VAL(11'b00000000000), .PCS_L64_R1_L64_BYPASS_TEST(1'b1)
        , .PCS_L64_R1_L64_CFG_TEST_PATTERN_EN(1'b0), .PCS_L64_R1_L64_CFG_TEST_PATT_TYPE_SEL(1'b0)
        , .PCS_L64_R1_L64_CFG_TEST_PRBS31_EN(1'b0), .PCS_L64_R1_L64_CFG_TEST_PATT_DATA_SEL(1'b0)
        , .PCS_L64_R2_L64_SEED_A_VALUE_LO32(32'b00000000000000000000000000000000)
        , .PCS_L64_R3_L64_SEED_A_VALUE_HI26(26'b00000000000000000000000000)
        , .PCS_L64_R4_L64_SEED_B_VALUE_LO32(32'b00000000000000000000000000000000)
        , .PCS_L64_R5_L64_SEED_B_VALUE_HI26(26'b00000000000000000000000000)
        , .PCS_L64_R6_L64_TX_ADV_CYC_DLY(5'b00000), .PCS_L64_R6_L64_TX_ADD_UI(16'b0000000000000000)
        , .PCS_L64_R7_L64_RX_ADV_CYC_DLY(5'b00000), .PCS_L64_R7_L64_RX_ADD_UI(16'b0000000000000000)
        , .PCS_L8_R0_L8_TXENCSWAPSEL(1'b0), .PCS_LRST_R0_LRST_SOFT_PCS_RX_RESET(1'b0)
        , .PCS_LRST_R0_LRST_SOFT_PCS_RX_DIV2_RESET(1'b0), .PCS_LRST_R0_LRST_ULCKD_CDR_RESETS_PCS_RX(1'b1)
        , .PCS_LRST_R0_LRST_SOFT_RXFWF_RESET(1'b0), .PCS_LRST_R0_LRST_SOFT_PCS_TX_RESET(1'b0)
        , .PCS_LRST_R0_LRST_SOFT_PCS_TX_DIV2_RESET(1'b0), .PCS_LRST_R0_LRST_ULCKD_PLL_RESETS_PCS_TX(1'b0)
        , .PCS_LRST_R0_LRST_SOFT_TXFWF_RESET(1'b0), .PCS_LRST_R0_LRST_SOFT_PIPE_RESET(7'b0000000)
        , .PCS_LRST_OPT_LRST_DISABLE_FAB_PCS_RESET_FOR_RX(1'b0), .PCS_LRST_OPT_LRST_DISABLE_FAB_PCS_RESET_FOR_TX(1'b0)
        , .PCS_OOB_R0_OOB_BURST_MIN_CYCLE(8'b00001111), .PCS_OOB_R0_OOB_BURST_MAX_CYCLE(8'b00010001)
        , .PCS_OOB_R0_OOB_WAKE_MIN_CYCLE(8'b00001111), .PCS_OOB_R0_OOB_WAKE_MAX_CYCLE(8'b00010001)
        , .PCS_OOB_R1_OOB_RST_INIT_MIN_CYCLE(8'b00101101), .PCS_OOB_R1_OOB_RST_INIT_MAX_CYCLE(8'b00110011)
        , .PCS_OOB_R1_OOB_SAS_MIN_CYCLE(8'b10001000), .PCS_OOB_R1_OOB_SAS_MAX_CYCLE(8'b10011000)
        , .PCS_OOB_R2_TXOOB_PROG_DATA_L32B(32'b00000000000000000000000000000000)
        , .PCS_OOB_R3_TXOOB_PROG_DATA_H8B(8'b00000000), .PCS_PMA_CTRL_R0_PMA_P2_ENTER_INT_MASK(1'b1)
        , .PCS_PMA_CTRL_R0_PMA_P2_EXIT_INT_MASK(1'b1), .PCS_PMA_CTRL_R0_PMA_P2_ENTER_INT(1'b0)
        , .PCS_PMA_CTRL_R0_PMA_P2_EXIT_INT(1'b0), .PCS_PMA_CTRL_R0_PMA_RXPLL_LOCK_INT_MASK(1'b1)
        , .PCS_PMA_CTRL_R0_PMA_RXPLL_UNLOCK_INT_MASK(1'b1), .PCS_PMA_CTRL_R0_PMA_RXPLL_LOCK_INT(1'b0)
        , .PCS_PMA_CTRL_R0_PMA_RXPLL_UNLOCK_INT(1'b0), .PCS_PMA_CTRL_R0_PMA_RXPLL_FLOCK_SEL(1'b0)
        , .PCS_PMA_CTRL_R0_PMA_TXPLL_LOCK_INT_MASK(1'b1), .PCS_PMA_CTRL_R0_PMA_TXPLL_UNLOCK_INT_MASK(1'b1)
        , .PCS_PMA_CTRL_R0_PMA_TXPLL_LOCK_INT(1'b0), .PCS_PMA_CTRL_R0_PMA_TXPLL_UNLOCK_INT(1'b0)
        , .PCS_PMA_CTRL_R1_RXBEACON_MAX_PULSE_WIDTH(11'b11001000000), .PCS_PMA_CTRL_R1_TXBEACON_PULSE_WIDTH(12'b000000001010)
        , .PCS_PMA_CTRL_R2_PD_PLL_CNT(8'b10100110), .PCS_PMA_CTRL_R2_PIPE_RATE_INIT(2'b00)
        , .PCS_PMA_CTRL_R2_FAB_DRIVES_TXPADS(1'b0), .PCS_MSTR_CTRL_LANE_MSTR(2'b00)
        , .MAIN_SOFT_RESET_PERIPH(1'b0), .MAIN_SOFT_RESET_NV_MAP(1'b0)
        , .MAIN_SOFT_RESET_V_MAP(1'b0), .MAIN_MAJOR_PCIE_USAGE_MODE(4'b1000)
        , .MAIN_INT_PIPE_CLK_CTRL_PCLK_INT_LN0_SEL(2'b10), .MAIN_INT_PIPE_CLK_CTRL_PCLK_INT_LN1_SEL(2'b10)
        , .MAIN_INT_PIPE_CLK_CTRL_PCLK_INT_LN2_SEL(1'b0), .MAIN_INT_PIPE_CLK_CTRL_PCLK_INT_LN3_SEL(1'b1)
        , .MAIN_EXT_PIPE_CLK_CTRL_PCLK_EXT_LN0_SEL(1'b0), .MAIN_EXT_PIPE_CLK_CTRL_PCLK_EXT_LN1_SEL(1'b0)
        , .MAIN_EXT_PIPE_CLK_CTRL_PCLK_EXT_LN2_SEL(1'b0), .MAIN_EXT_PIPE_CLK_CTRL_PCLK_EXT_LN3_SEL(1'b0)
        , .MAIN_QMUX_R0_PCIE_DBG_SEL(3'b111), .MAIN_DLL_CTRL0_PHASE_P(2'b11)
        , .MAIN_DLL_CTRL0_PHASE_S(2'b11), .MAIN_DLL_CTRL0_SEL_P(2'b00)
        , .MAIN_DLL_CTRL0_SEL_S(2'b00), .MAIN_DLL_CTRL0_REF_SEL(1'b0)
        , .MAIN_DLL_CTRL0_FB_SEL(1'b0), .MAIN_DLL_CTRL0_DIV_SEL(1'b0)
        , .MAIN_DLL_CTRL0_ALU_UPD(2'b00), .MAIN_DLL_CTRL0_LOCK_FRC(1'b0)
        , .MAIN_DLL_CTRL0_LOCK_FLT(2'b00), .MAIN_DLL_CTRL0_LOCK_HIGH(4'b1000)
        , .MAIN_DLL_CTRL0_LOCK_LOW(4'b1000), .MAIN_DLL_CTRL1_SET_ALU(8'b00000000)
        , .MAIN_DLL_CTRL1_ADJ_DEL4(7'b0000000), .MAIN_DLL_CTRL1_TEST_S(1'b0)
        , .MAIN_DLL_CTRL1_TEST_RING(1'b0), .MAIN_DLL_CTRL1_INIT_CODE(6'b000000)
        , .MAIN_DLL_CTRL1_RELOCK_FAST(1'b0), .MAIN_DLL_STAT0_RESET(1'b0)
        , .MAIN_DLL_STAT0_PHASE_MOVE_CLK(1'b0), .MAIN_OVRLY_AXI0_IFC_MODE(2'b01)
        , .MAIN_OVRLY_AXI1_IFC_MODE(2'b01), .MAIN_INT_PIPE_CLK_CTRL_PCIE_0_PCLK_SEL(3'b110)
        , .MAIN_INT_PIPE_CLK_CTRL_PCIE_1_PCLK_SEL(3'b010), .MAIN_CLK_CTRL_AXI0_CLKENA(1'b0)
        , .MAIN_CLK_CTRL_AXI1_CLKENA(1'b0), .MAIN_DLL_STAT0_LOCK_INT_EN(1'b0)
        , .MAIN_DLL_STAT0_UNLOCK_INT_EN(1'b0), .MAIN_DLL_STAT0_LOCK_INT(1'b0)
        , .MAIN_DLL_STAT0_UNLOCK_INT(1'b1), .MAIN_TEST_DLL_RING_OSC_ENABLE(1'b0)
        , .MAIN_TEST_DLL_REF_ENABLE(1'b0), .MAIN_SPARE_SCRATCHPAD(8'b00000000)
        , .MAIN_SPARE_SPARE_CTRL(24'b000000000000000000000000), .PMA_SOFT_RESET_PERIPH(1'b0)
        , .PMA_DES_CDR_CTRL_3_CST1_CDR(2'b00), .PMA_DES_CDR_CTRL_3_CST2_CDR(2'b00)
        , .PMA_DES_CDR_CTRL_3_RST1_CDR(2'b00), .PMA_DES_CDR_CTRL_3_RST2_CDR(2'b00)
        , .PMA_DES_CDR_CTRL_3_RXDRV_CDR(2'b00), .PMA_DES_DFEEM_CTRL_3_CST1_DFEEM(2'b00)
        , .PMA_DES_DFEEM_CTRL_3_CST2_DFEEM(2'b00), .PMA_DES_DFEEM_CTRL_3_RST1_DFEEM(2'b00)
        , .PMA_DES_DFEEM_CTRL_3_RST2_DFEEM(2'b00), .PMA_DES_DFE_CTRL_2_RXDRV_DFE(2'b00)
        , .PMA_DES_DFE_CTRL_2_CTLEEN_DFE(1'b0), .PMA_DES_EM_CTRL_2_RXDRV_EM(2'b00)
        , .PMA_DES_EM_CTRL_2_CTLEEN_EM(1'b0), .PMA_DES_IN_TERM_RXRTRIM(4'b0111)
        , .PMA_DES_IN_TERM_RXTEN(1'b0), .PMA_DES_IN_TERM_RXRTRIM_SEL(2'b01)
        , .PMA_DES_IN_TERM_ACCOUPLE_RXVCM_EN(1'b1), .PMA_DES_PKDET_RXPKDETEN(1'b1)
        , .PMA_DES_PKDET_RXPKDETRANGE(1'b0), .PMA_DES_PKDET_RXPKDET_LOW_THRESHOLD(3'b001)
        , .PMA_DES_PKDET_RXPKDET_HIGH_THRESHOLD(3'b010), .PMA_DES_RTL_LOCK_CTRL_LOCK_MODE(1'b0)
        , .PMA_DES_RTL_LOCK_CTRL_LOCK_OVERRIDE(2'b00), .PMA_DES_RTL_LOCK_CTRL_FDET_SAMPLE_PERIODS(5'b00001)
        , .PMA_DES_RXPLL_DIV_RXPLL_FBDIV(8'b00110010), .PMA_DES_RXPLL_DIV_RXPLL_REFDIV(5'b00010)
        , .PMA_DES_RXPLL_DIV_RXPLL_RANGE(2'b00), .PMA_DES_RXPLL_DIV_CDR_GAIN(1'b0)
        , .PMA_DES_TEST_BUS_RXATESTEN(1'b0), .PMA_DES_CLK_CTRL_RXREFCLK_SEL(3'b100)
        , .PMA_DES_CLK_CTRL_DESMODE(3'b111), .PMA_DES_CLK_CTRL_DATALOCKEN(1'b0)
        , .PMA_DES_CLK_CTRL_DATALOCKDIVEN(1'b0), .PMA_SER_CTRL_TXVBGREF_SEL(1'b0)
        , .PMA_SER_CLK_CTRL_TXPOSTDIVEN(1'b0), .PMA_SER_CLK_CTRL_TXPOSTDIV(2'b00)
        , .PMA_SER_CLK_CTRL_TXBITCLKSEL(1'b0), .PMA_SER_CLK_CTRL_SERMODE(3'b111)
        , .PMA_SER_DRV_BYP_BYPASS_VALUE(8'b00000000), .PMA_SER_DRV_BYP_TX_BYPASS_SELECT_RTL(2'b00)
        , .PMA_SER_DRV_BYP_TX_BYPASS_SELECT(1'b0), .PMA_SER_RXDET_CTRL_RXDETECT_STEP_WAIT_COUNT(5'b10000)
        , .PMA_SER_TERM_CTRL_TXCM_LEVEL(2'b00), .PMA_SER_TERM_CTRL_TXTEN(1'b0)
        , .PMA_SER_TERM_CTRL_TXRTRIM_SEL(2'b01), .PMA_SER_TERM_CTRL_TXRTRIM(4'b0111)
        , .PMA_SER_TEST_BUS_TXATESTEN(1'b0), .PMA_SER_DRV_DATA_CTRL_TXDEL(16'b0000000000000000)
        , .PMA_SER_DRV_DATA_CTRL_TXDATA_INV(8'b00000000), .PMA_SER_DRV_CTRL_TXDRVTRIM(24'b000000000000000000000000)
        , .PMA_SER_DRV_CTRL_TXDRV(3'b001), .PMA_SER_DRV_CTRL_TXITRIM(2'b10)
        , .PMA_SER_DRV_CTRL_TXODRV(2'b00), .PMA_SER_DRV_CTRL_SEL_TXDRV_CTRL_SEL(1'b0)
        , .PMA_SER_DRV_CTRL_SEL_TXODRV_BOOSTER(1'b0), .PMA_SER_DRV_CTRL_SEL_TXMARGIN(3'b000)
        , .PMA_SER_DRV_CTRL_SEL_TXSWING(1'b0), .PMA_SER_DRV_CTRL_SEL_TXDEEMPHASIS(1'b0)
        , .PMA_SER_DRV_CTRL_SEL_TXDEEMPHASIS_BEACON(1'b0), .PMA_SERDES_RTL_CTRL_RX_HALF_RATE10BIT(1'b0)
        , .PMA_SERDES_RTL_CTRL_TX_HALF_RATE10BIT(1'b0), .PCS_SOFT_RESET_PERIPH(1'b0)
        , .PCS_LFWF_R0_RXFWF_RATIO(2'b00), .PCS_LFWF_R0_TXFWF_RATIO(2'b00)
        , .PCS_LOVR_R0_FAB_IFC_MODE(4'b0000), .PCS_LOVR_R0_PCSPMA_IFC_MODE(4'b0001)
        , .PCS_LPIP_R0_PIPEENABLE(1'b1), .PCS_LPIP_R0_PIPEMODE(1'b0), .PCS_LPIP_R0_PIPE_PCIE_HC(1'b1)
        , .PCS_L64_R0_L64_CFG_BYPASS_SCRAMBLER(1'b0), .PCS_L64_R0_L64_CFG_BYPASS_DISPARITY(1'b1)
        , .PCS_L64_R0_L64_CFG_BYPASS_GEARBOX(1'b0), .PCS_L64_R0_L64_CFG_GRBX_64B67B(1'b0)
        , .PCS_L64_R0_L64_CFG_BER_MON_EN(1'b1), .PCS_L64_R0_L64_CFG_BYPASS_8B_MODE(1'b0)
        , .PCS_L64_R0_L64_CFG_GRBX_SM_C49(1'b0), .PCS_L64_R0_L64_CFG_GRBX_SM_C82(1'b0)
        , .PCS_L8_R0_L8_GEARMODE(2'b00), .PCS_LNTV_R0_LNTV_RX_GEAR(1'b0)
        , .PCS_LNTV_R0_LNTV_RX_IN_WIDTH(3'b111), .PCS_LNTV_R0_LNTV_RX_MODE(1'b0)
        , .PCS_LNTV_R0_LNTV_TX_GEAR(1'b0), .PCS_LNTV_R0_LNTV_TX_OUT_WIDTH(3'b111)
        , .PCS_LNTV_R0_LNTV_TX_MODE(1'b0), .PCS_LCLK_R0_LCLK_EPCS_RX_CLK_SEL(2'b00)
        , .PCS_LCLK_R0_LCLK_EPCS_TX_CLK_SEL(2'b00), .PCS_LCLK_R0_LCLK_TXFWF_TMG_MODE(1'b0)
        , .PCS_LCLK_R0_LCLK_PCS_RX_CLK_SEL(2'b11), .PCS_LCLK_R0_LCLK_PCS_TX_CLK_SEL(2'b11)
        , .PCS_LCLK_R0_LCLK_RXFWF_WCLK_SEL(2'b00), .PCS_LCLK_R0_LCLK_TXFWF_RCLK_SEL(2'b00)
        , .PCS_LCLK_R0_LCLK_RXFWF_WCLK_PIPE(1'b0), .PCS_LCLK_R1_LCLK_ENA_64B6XB_RX_CLK(1'b0)
        , .PCS_LCLK_R1_LCLK_ENA_64B6XB_RX_CLK_DIV2(1'b0), .PCS_LCLK_R1_LCLK_ENA_64B6XB_TX_CLK(1'b0)
        , .PCS_LCLK_R1_LCLK_ENA_64B6XB_TX_CLK_DIV2(1'b0), .PCS_LCLK_R1_LCLK_ENA_8B10B_RX_CLK(1'b0)
        , .PCS_LCLK_R1_LCLK_ENA_8B10B_RXFWF_WCLK(1'b0), .PCS_LCLK_R1_LCLK_ENA_8B10B_TX_CLK(1'b0)
        , .PCS_LCLK_R1_LCLK_ENA_8B10B_TXFWF_RCLK(1'b0), .PCS_LCLK_R1_LCLK_ENA_NATIVE_RX_CLK(1'b0)
        , .PCS_LCLK_R1_LCLK_ENA_NATIVE_RXFWF_WCLK(1'b0), .PCS_LCLK_R1_LCLK_ENA_NATIVE_TX_CLK(1'b0)
        , .PCS_LCLK_R1_LCLK_ENA_NATIVE_TXFWF_RCLK(1'b0), .PCS_LCLK_R1_LCLK_ENA_PIPE_LCL(1'b1)
        , .PCS_LCLK_R1_LCLK_ENA_PIPE_OUT(1'b1), .PCS_PMA_CTRL_R0_PIPE_P0S_EN(1'b1)
        , .PCS_PMA_CTRL_R0_PIPE_P1_EN(1'b1), .PCS_PMA_CTRL_R0_PIPE_P2_EN(1'b1)
        , .PCS_PMA_CTRL_R0_FLASH_FREEZE_P0S_EN(1'b0), .PCS_PMA_CTRL_R0_FLASH_FREEZE_P1_EN(1'b0)
        , .PCS_PMA_CTRL_R0_FLASH_FREEZE_P2_EN(1'b0), .PCS_PMA_CTRL_R0_FAB_EPCS_PMA_RESET_B_EN(1'b1)
         )  PCIESS_LANE2_Pipe_AXI1 (.M_ARADDR_31(
        PCIESS_AXI_1_M_ARADDR[31]), .M_ARADDR_30(
        PCIESS_AXI_1_M_ARADDR[30]), .M_ARADDR_29(
        PCIESS_AXI_1_M_ARADDR[29]), .M_ARADDR_28(
        PCIESS_AXI_1_M_ARADDR[28]), .M_ARADDR_0(
        PCIESS_AXI_1_M_ARADDR[0]), .M_ARADDR_1(
        PCIESS_AXI_1_M_ARADDR[1]), .M_ARADDR_2(
        PCIESS_AXI_1_M_ARADDR[2]), .M_ARADDR_3(
        PCIESS_AXI_1_M_ARADDR[3]), .M_ARADDR_4(
        PCIESS_AXI_1_M_ARADDR[4]), .M_ARADDR_5(
        PCIESS_AXI_1_M_ARADDR[5]), .M_ARADDR_6(
        PCIESS_AXI_1_M_ARADDR[6]), .M_ARADDR_7(
        PCIESS_AXI_1_M_ARADDR[7]), .M_ARADDR_8(
        PCIESS_AXI_1_M_ARADDR[8]), .M_ARADDR_9(
        PCIESS_AXI_1_M_ARADDR[9]), .M_ARADDR_10(
        PCIESS_AXI_1_M_ARADDR[10]), .M_ARADDR_11(
        PCIESS_AXI_1_M_ARADDR[11]), .M_ARADDR_12(
        PCIESS_AXI_1_M_ARADDR[12]), .M_ARADDR_13(
        PCIESS_AXI_1_M_ARADDR[13]), .M_ARADDR_14(
        PCIESS_AXI_1_M_ARADDR[14]), .M_ARADDR_15(
        PCIESS_AXI_1_M_ARADDR[15]), .M_ARADDR_16(
        PCIESS_AXI_1_M_ARADDR[16]), .M_ARADDR_17(
        PCIESS_AXI_1_M_ARADDR[17]), .M_ARADDR_18(
        PCIESS_AXI_1_M_ARADDR[18]), .M_ARADDR_19(
        PCIESS_AXI_1_M_ARADDR[19]), .M_ARADDR_20(
        PCIESS_AXI_1_M_ARADDR[20]), .M_ARADDR_21(
        PCIESS_AXI_1_M_ARADDR[21]), .M_ARADDR_22(
        PCIESS_AXI_1_M_ARADDR[22]), .M_ARADDR_23(
        PCIESS_AXI_1_M_ARADDR[23]), .S_RDATA({PCIESS_AXI_1_S_RDATA[63], 
        PCIESS_AXI_1_S_RDATA[62], PCIESS_AXI_1_S_RDATA[61], 
        PCIESS_AXI_1_S_RDATA[60], PCIESS_AXI_1_S_RDATA[59], 
        PCIESS_AXI_1_S_RDATA[58], PCIESS_AXI_1_S_RDATA[57], 
        PCIESS_AXI_1_S_RDATA[56], PCIESS_AXI_1_S_RDATA[55], 
        PCIESS_AXI_1_S_RDATA[54], PCIESS_AXI_1_S_RDATA[53], 
        PCIESS_AXI_1_S_RDATA[52], PCIESS_AXI_1_S_RDATA[51], 
        PCIESS_AXI_1_S_RDATA[50], PCIESS_AXI_1_S_RDATA[49], 
        PCIESS_AXI_1_S_RDATA[48], PCIESS_AXI_1_S_RDATA[47], 
        PCIESS_AXI_1_S_RDATA[46], PCIESS_AXI_1_S_RDATA[45], 
        PCIESS_AXI_1_S_RDATA[44], PCIESS_AXI_1_S_RDATA[43], 
        PCIESS_AXI_1_S_RDATA[42], PCIESS_AXI_1_S_RDATA[41], 
        PCIESS_AXI_1_S_RDATA[40], PCIESS_AXI_1_S_RDATA[39], 
        PCIESS_AXI_1_S_RDATA[38], PCIESS_AXI_1_S_RDATA[37], 
        PCIESS_AXI_1_S_RDATA[36], PCIESS_AXI_1_S_RDATA[35], 
        PCIESS_AXI_1_S_RDATA[34], PCIESS_AXI_1_S_RDATA[33], 
        PCIESS_AXI_1_S_RDATA[32], PCIESS_AXI_1_S_RDATA[31], 
        PCIESS_AXI_1_S_RDATA[30], PCIESS_AXI_1_S_RDATA[29], 
        PCIESS_AXI_1_S_RDATA[28], PCIESS_AXI_1_S_RDATA[27], 
        PCIESS_AXI_1_S_RDATA[26], PCIESS_AXI_1_S_RDATA[25], 
        PCIESS_AXI_1_S_RDATA[24], PCIESS_AXI_1_S_RDATA[23], 
        PCIESS_AXI_1_S_RDATA[22], PCIESS_AXI_1_S_RDATA[21], 
        PCIESS_AXI_1_S_RDATA[20], PCIESS_AXI_1_S_RDATA[19], 
        PCIESS_AXI_1_S_RDATA[18], PCIESS_AXI_1_S_RDATA[17], 
        PCIESS_AXI_1_S_RDATA[16], PCIESS_AXI_1_S_RDATA[15], 
        PCIESS_AXI_1_S_RDATA[14], PCIESS_AXI_1_S_RDATA[13], 
        PCIESS_AXI_1_S_RDATA[12], PCIESS_AXI_1_S_RDATA[11], 
        PCIESS_AXI_1_S_RDATA[10], PCIESS_AXI_1_S_RDATA[9], 
        PCIESS_AXI_1_S_RDATA[8], PCIESS_AXI_1_S_RDATA[7], 
        PCIESS_AXI_1_S_RDATA[6], PCIESS_AXI_1_S_RDATA[5], 
        PCIESS_AXI_1_S_RDATA[4], PCIESS_AXI_1_S_RDATA[3], 
        PCIESS_AXI_1_S_RDATA[2], PCIESS_AXI_1_S_RDATA[1], 
        PCIESS_AXI_1_S_RDATA[0]}), .RX_REF_CLK(gnd_net), .S_ARADDR_31(
        PCIESS_AXI_1_S_ARADDR[31]), .S_ARADDR_30(
        PCIESS_AXI_1_S_ARADDR[30]), .S_ARADDR_28(
        PCIESS_AXI_1_S_ARADDR[28]), .S_ARADDR_0(
        PCIESS_AXI_1_S_ARADDR[0]), .S_ARADDR_1(
        PCIESS_AXI_1_S_ARADDR[1]), .S_ARADDR_2(
        PCIESS_AXI_1_S_ARADDR[2]), .S_ARADDR_3(
        PCIESS_AXI_1_S_ARADDR[3]), .S_ARADDR_4(
        PCIESS_AXI_1_S_ARADDR[4]), .S_ARADDR_5(
        PCIESS_AXI_1_S_ARADDR[5]), .S_ARADDR_6(
        PCIESS_AXI_1_S_ARADDR[6]), .S_ARADDR_7(
        PCIESS_AXI_1_S_ARADDR[7]), .S_ARADDR_8(
        PCIESS_AXI_1_S_ARADDR[8]), .S_ARADDR_9(
        PCIESS_AXI_1_S_ARADDR[9]), .S_ARADDR_10(
        PCIESS_AXI_1_S_ARADDR[10]), .S_ARADDR_11(
        PCIESS_AXI_1_S_ARADDR[11]), .S_ARADDR_12(
        PCIESS_AXI_1_S_ARADDR[12]), .S_ARADDR_13(
        PCIESS_AXI_1_S_ARADDR[13]), .S_ARADDR_14(
        PCIESS_AXI_1_S_ARADDR[14]), .S_ARADDR_15(
        PCIESS_AXI_1_S_ARADDR[15]), .S_ARADDR_16(
        PCIESS_AXI_1_S_ARADDR[16]), .S_ARADDR_17(
        PCIESS_AXI_1_S_ARADDR[17]), .S_ARADDR_18(
        PCIESS_AXI_1_S_ARADDR[18]), .S_ARADDR_19(
        PCIESS_AXI_1_S_ARADDR[19]), .S_ARADDR_20(
        PCIESS_AXI_1_S_ARADDR[20]), .S_ARADDR_21(
        PCIESS_AXI_1_S_ARADDR[21]), .S_ARADDR_22(
        PCIESS_AXI_1_S_ARADDR[22]), .S_ARADDR_23(
        PCIESS_AXI_1_S_ARADDR[23]), .S_WDATA({PCIESS_AXI_1_S_WDATA[63], 
        PCIESS_AXI_1_S_WDATA[62], PCIESS_AXI_1_S_WDATA[61], 
        PCIESS_AXI_1_S_WDATA[60], PCIESS_AXI_1_S_WDATA[59], 
        PCIESS_AXI_1_S_WDATA[58], PCIESS_AXI_1_S_WDATA[57], 
        PCIESS_AXI_1_S_WDATA[56], PCIESS_AXI_1_S_WDATA[55], 
        PCIESS_AXI_1_S_WDATA[54], PCIESS_AXI_1_S_WDATA[53], 
        PCIESS_AXI_1_S_WDATA[52], PCIESS_AXI_1_S_WDATA[51], 
        PCIESS_AXI_1_S_WDATA[50], PCIESS_AXI_1_S_WDATA[49], 
        PCIESS_AXI_1_S_WDATA[48], PCIESS_AXI_1_S_WDATA[47], 
        PCIESS_AXI_1_S_WDATA[46], PCIESS_AXI_1_S_WDATA[45], 
        PCIESS_AXI_1_S_WDATA[44], PCIESS_AXI_1_S_WDATA[43], 
        PCIESS_AXI_1_S_WDATA[42], PCIESS_AXI_1_S_WDATA[41], 
        PCIESS_AXI_1_S_WDATA[40], PCIESS_AXI_1_S_WDATA[39], 
        PCIESS_AXI_1_S_WDATA[38], PCIESS_AXI_1_S_WDATA[37], 
        PCIESS_AXI_1_S_WDATA[36], PCIESS_AXI_1_S_WDATA[35], 
        PCIESS_AXI_1_S_WDATA[34], PCIESS_AXI_1_S_WDATA[33], 
        PCIESS_AXI_1_S_WDATA[32], PCIESS_AXI_1_S_WDATA[31], 
        PCIESS_AXI_1_S_WDATA[30], PCIESS_AXI_1_S_WDATA[29], 
        PCIESS_AXI_1_S_WDATA[28], PCIESS_AXI_1_S_WDATA[27], 
        PCIESS_AXI_1_S_WDATA[26], PCIESS_AXI_1_S_WDATA[25], 
        PCIESS_AXI_1_S_WDATA[24], PCIESS_AXI_1_S_WDATA[23], 
        PCIESS_AXI_1_S_WDATA[22], PCIESS_AXI_1_S_WDATA[21], 
        PCIESS_AXI_1_S_WDATA[20], PCIESS_AXI_1_S_WDATA[19], 
        PCIESS_AXI_1_S_WDATA[18], PCIESS_AXI_1_S_WDATA[17], 
        PCIESS_AXI_1_S_WDATA[16], PCIESS_AXI_1_S_WDATA[15], 
        PCIESS_AXI_1_S_WDATA[14], PCIESS_AXI_1_S_WDATA[13], 
        PCIESS_AXI_1_S_WDATA[12], PCIESS_AXI_1_S_WDATA[11], 
        PCIESS_AXI_1_S_WDATA[10], PCIESS_AXI_1_S_WDATA[9], 
        PCIESS_AXI_1_S_WDATA[8], PCIESS_AXI_1_S_WDATA[7], 
        PCIESS_AXI_1_S_WDATA[6], PCIESS_AXI_1_S_WDATA[5], 
        PCIESS_AXI_1_S_WDATA[4], PCIESS_AXI_1_S_WDATA[3], 
        PCIESS_AXI_1_S_WDATA[2], PCIESS_AXI_1_S_WDATA[1], 
        PCIESS_AXI_1_S_WDATA[0]}), .M_ARADDR_HW_0(
        PCIE_1_M_ARADDR_0_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_0_net), 
        .M_ARADDR_HW_1(
        PCIE_1_M_ARADDR_1_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_1_net), 
        .M_ARADDR_HW_2(
        PCIE_1_M_ARADDR_2_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_2_net), 
        .M_ARADDR_HW_3(
        PCIE_1_M_ARADDR_3_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_3_net), 
        .M_ARADDR_HW_4(
        PCIE_1_M_ARADDR_4_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_4_net), 
        .M_ARADDR_HW_5(
        PCIE_1_M_ARADDR_5_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_5_net), 
        .M_ARADDR_HW_6(
        PCIE_1_M_ARADDR_6_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_6_net), 
        .M_ARADDR_HW_7(
        PCIE_1_M_ARADDR_7_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_7_net), 
        .M_ARADDR_HW_8(
        PCIE_1_M_ARADDR_8_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_8_net), 
        .M_ARADDR_HW_9(
        PCIE_1_M_ARADDR_9_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_9_net), 
        .M_ARADDR_HW_10(
        PCIE_1_M_ARADDR_10_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_10_net), 
        .M_ARADDR_HW_11(
        PCIE_1_M_ARADDR_11_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_11_net), 
        .M_ARADDR_HW_12(
        PCIE_1_M_ARADDR_12_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_12_net), 
        .M_ARADDR_HW_13(
        PCIE_1_M_ARADDR_13_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_13_net), 
        .M_ARADDR_HW_14(
        PCIE_1_M_ARADDR_14_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_14_net), 
        .M_ARADDR_HW_15(
        PCIE_1_M_ARADDR_15_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_15_net), 
        .M_ARADDR_HW_16(
        PCIE_1_M_ARADDR_16_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_16_net), 
        .M_ARADDR_HW_17(
        PCIE_1_M_ARADDR_17_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_17_net), 
        .M_ARADDR_HW_18(
        PCIE_1_M_ARADDR_18_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_18_net), 
        .M_ARADDR_HW_19(
        PCIE_1_M_ARADDR_19_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_19_net), 
        .M_ARADDR_HW_20(
        PCIE_1_M_ARADDR_20_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_20_net), 
        .M_ARADDR_HW_21(
        PCIE_1_M_ARADDR_21_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_21_net), 
        .M_ARADDR_HW_22(
        PCIE_1_M_ARADDR_22_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_22_net), 
        .M_ARADDR_HW_23(
        PCIE_1_M_ARADDR_23_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_23_net), 
        .M_ARADDR_HW_28(
        PCIE_1_M_ARADDR_28_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_28_net), 
        .M_ARADDR_HW_29(
        PCIE_1_M_ARADDR_29_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_29_net), 
        .M_ARADDR_HW_30(
        PCIE_1_M_ARADDR_30_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_30_net), 
        .M_ARADDR_HW_31(
        PCIE_1_M_ARADDR_31_PCIESS_LANE2_Pipe_AXI1_M_ARADDR_HW_31_net), 
        .S_ARADDR_HW_0(
        PCIE_1_S_ARADDR_0_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_0_net), 
        .S_ARADDR_HW_1(
        PCIE_1_S_ARADDR_1_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_1_net), 
        .S_ARADDR_HW_2(
        PCIE_1_S_ARADDR_2_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_2_net), 
        .S_ARADDR_HW_3(
        PCIE_1_S_ARADDR_3_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_3_net), 
        .S_ARADDR_HW_4(
        PCIE_1_S_ARADDR_4_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_4_net), 
        .S_ARADDR_HW_5(
        PCIE_1_S_ARADDR_5_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_5_net), 
        .S_ARADDR_HW_6(
        PCIE_1_S_ARADDR_6_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_6_net), 
        .S_ARADDR_HW_7(
        PCIE_1_S_ARADDR_7_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_7_net), 
        .S_ARADDR_HW_8(
        PCIE_1_S_ARADDR_8_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_8_net), 
        .S_ARADDR_HW_9(
        PCIE_1_S_ARADDR_9_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_9_net), 
        .S_ARADDR_HW_10(
        PCIE_1_S_ARADDR_10_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_10_net), 
        .S_ARADDR_HW_11(
        PCIE_1_S_ARADDR_11_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_11_net), 
        .S_ARADDR_HW_12(
        PCIE_1_S_ARADDR_12_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_12_net), 
        .S_ARADDR_HW_13(
        PCIE_1_S_ARADDR_13_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_13_net), 
        .S_ARADDR_HW_14(
        PCIE_1_S_ARADDR_14_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_14_net), 
        .S_ARADDR_HW_15(
        PCIE_1_S_ARADDR_15_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_15_net), 
        .S_ARADDR_HW_16(
        PCIE_1_S_ARADDR_16_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_16_net), 
        .S_ARADDR_HW_17(
        PCIE_1_S_ARADDR_17_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_17_net), 
        .S_ARADDR_HW_18(
        PCIE_1_S_ARADDR_18_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_18_net), 
        .S_ARADDR_HW_19(
        PCIE_1_S_ARADDR_19_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_19_net), 
        .S_ARADDR_HW_20(
        PCIE_1_S_ARADDR_20_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_20_net), 
        .S_ARADDR_HW_21(
        PCIE_1_S_ARADDR_21_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_21_net), 
        .S_ARADDR_HW_22(
        PCIE_1_S_ARADDR_22_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_22_net), 
        .S_ARADDR_HW_23(
        PCIE_1_S_ARADDR_23_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_23_net), 
        .S_ARADDR_HW_28(
        PCIE_1_S_ARADDR_28_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_28_net), 
        .S_ARADDR_HW_30(
        PCIE_1_S_ARADDR_30_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_30_net), 
        .S_ARADDR_HW_31(
        PCIE_1_S_ARADDR_31_PCIESS_LANE2_Pipe_AXI1_S_ARADDR_HW_31_net), 
        .S_RDATA_HW({
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_63, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_62, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_61, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_60, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_59, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_58, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_57, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_56, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_55, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_54, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_53, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_52, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_51, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_50, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_49, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_48, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_47, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_46, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_45, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_44, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_43, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_42, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_41, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_40, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_39, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_38, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_37, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_36, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_35, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_34, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_33, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_32, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_31, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_30, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_29, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_28, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_27, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_26, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_25, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_24, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_23, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_22, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_21, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_20, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_19, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_18, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_17, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_16, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_15, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_14, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_13, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_12, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_11, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_10, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_9, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_8, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_7, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_6, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_5, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_4, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_3, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_2, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_1, 
        PCIE_1_S_RDATA_PCIESS_LANE2_Pipe_AXI1_S_RDATA_HW_net_0}), 
        .S_WDATA_HW({
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_63, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_62, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_61, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_60, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_59, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_58, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_57, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_56, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_55, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_54, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_53, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_52, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_51, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_50, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_49, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_48, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_47, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_46, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_45, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_44, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_43, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_42, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_41, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_40, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_39, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_38, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_37, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_36, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_35, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_34, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_33, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_32, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_31, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_30, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_29, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_28, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_27, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_26, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_25, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_24, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_23, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_22, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_21, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_20, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_19, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_18, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_17, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_16, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_15, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_14, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_13, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_12, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_11, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_10, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_9, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_8, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_7, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_6, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_5, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_4, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_3, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_2, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_1, 
        PCIE_1_S_WDATA_PCIESS_LANE2_Pipe_AXI1_S_WDATA_HW_net_0}), 
        .PCS_DEBUG({
        PCIE_COMMON_INSTANCE_PCS_DEBUG_2_PCIESS_LANE2_Pipe_AXI1_PCS_DEBUG_net_19, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_2_PCIESS_LANE2_Pipe_AXI1_PCS_DEBUG_net_18, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_2_PCIESS_LANE2_Pipe_AXI1_PCS_DEBUG_net_17, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_2_PCIESS_LANE2_Pipe_AXI1_PCS_DEBUG_net_16, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_2_PCIESS_LANE2_Pipe_AXI1_PCS_DEBUG_net_15, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_2_PCIESS_LANE2_Pipe_AXI1_PCS_DEBUG_net_14, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_2_PCIESS_LANE2_Pipe_AXI1_PCS_DEBUG_net_13, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_2_PCIESS_LANE2_Pipe_AXI1_PCS_DEBUG_net_12, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_2_PCIESS_LANE2_Pipe_AXI1_PCS_DEBUG_net_11, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_2_PCIESS_LANE2_Pipe_AXI1_PCS_DEBUG_net_10, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_2_PCIESS_LANE2_Pipe_AXI1_PCS_DEBUG_net_9, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_2_PCIESS_LANE2_Pipe_AXI1_PCS_DEBUG_net_8, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_2_PCIESS_LANE2_Pipe_AXI1_PCS_DEBUG_net_7, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_2_PCIESS_LANE2_Pipe_AXI1_PCS_DEBUG_net_6, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_2_PCIESS_LANE2_Pipe_AXI1_PCS_DEBUG_net_5, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_2_PCIESS_LANE2_Pipe_AXI1_PCS_DEBUG_net_4, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_2_PCIESS_LANE2_Pipe_AXI1_PCS_DEBUG_net_3, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_2_PCIESS_LANE2_Pipe_AXI1_PCS_DEBUG_net_2, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_2_PCIESS_LANE2_Pipe_AXI1_PCS_DEBUG_net_1, 
        PCIE_COMMON_INSTANCE_PCS_DEBUG_2_PCIESS_LANE2_Pipe_AXI1_PCS_DEBUG_net_0})
        , .REF_CLK_N(gnd_net), .REF_CLK_P(PCIESS_LANE2_CDR_REF_CLK_0), 
        .RX_N(PCIESS_LANE_RXD2_N), .RX_P(PCIESS_LANE_RXD2_P), .TX_N(
        PCIESS_LANE_TXD2_N), .TX_P(PCIESS_LANE_TXD2_P), .JA_CLK(), 
        .TX_BIT_CLK_0(PCIE_1_TX_BIT_CLK), .TX_BIT_CLK_1(gnd_net), 
        .TX_PLL_LOCK_0(PCIE_1_TX_PLL_LOCK), .TX_PLL_LOCK_1(gnd_net), 
        .TX_PLL_REF_CLK_0(PCIE_1_TX_PLL_REF_CLK), .TX_PLL_REF_CLK_1(
        gnd_net), .TX_CLK_G(), .RX_CLK_G(), .PMA_DEBUG(
        PCIE_COMMON_INSTANCE_PMA_DEBUG_2_PCIESS_LANE2_Pipe_AXI1_PMA_DEBUG_net)
        , .ARST_N({nc345, nc346}), .DRI_CLK(gnd_net), .DRI_CTRL({
        gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, 
        gnd_net, gnd_net, gnd_net, gnd_net}), .DRI_WDATA({gnd_net, 
        gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, 
        gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, 
        gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, 
        gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, gnd_net, 
        gnd_net, gnd_net, gnd_net, gnd_net}), .DRI_ARST_N(vcc_net), 
        .DRI_RDATA({nc347, nc348, nc349, nc350, nc351, nc352, nc353, 
        nc354, nc355, nc356, nc357, nc358, nc359, nc360, nc361, nc362, 
        nc363, nc364, nc365, nc366, nc367, nc368, nc369, nc370, nc371, 
        nc372, nc373, nc374, nc375, nc376, nc377, nc378, nc379}), 
        .DRI_INTERRUPT(), .PHYSTATUS_0(
        PCIE_1_PHYSTATUS_2_PCIESS_LANE2_Pipe_AXI1_PHYSTATUS_0_net), 
        .POWERDOWN({
        PCIE_1_POWERDOWN_PCIESS_LANE2_Pipe_AXI1_POWERDOWN_net_1, 
        PCIE_1_POWERDOWN_PCIESS_LANE2_Pipe_AXI1_POWERDOWN_net_0}), 
        .RATE({PCIE_1_RATE_PCIESS_LANE2_Pipe_AXI1_RATE_net_1, 
        PCIE_1_RATE_PCIESS_LANE2_Pipe_AXI1_RATE_net_0}), .RESET_N(
        PCIE_1_RESET_N_PCIESS_LANE2_Pipe_AXI1_RESET_N_net), .RXDATA_0({
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_31, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_30, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_29, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_28, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_27, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_26, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_25, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_24, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_23, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_22, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_21, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_20, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_19, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_18, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_17, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_16, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_15, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_14, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_13, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_12, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_11, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_10, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_9, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_8, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_7, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_6, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_5, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_4, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_3, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_2, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_1, 
        PCIE_1_RXDATA_2_PCIESS_LANE2_Pipe_AXI1_RXDATA_0_net_0}), 
        .RXDATAK_0({
        PCIE_1_RXDATAK_2_PCIESS_LANE2_Pipe_AXI1_RXDATAK_0_net_3, 
        PCIE_1_RXDATAK_2_PCIESS_LANE2_Pipe_AXI1_RXDATAK_0_net_2, 
        PCIE_1_RXDATAK_2_PCIESS_LANE2_Pipe_AXI1_RXDATAK_0_net_1, 
        PCIE_1_RXDATAK_2_PCIESS_LANE2_Pipe_AXI1_RXDATAK_0_net_0}), 
        .RXELECIDLE_0(
        PCIE_1_RXELECIDLE_2_PCIESS_LANE2_Pipe_AXI1_RXELECIDLE_0_net), 
        .RXPOLARITY_0(
        PCIE_1_RXPOLARITY_2_PCIESS_LANE2_Pipe_AXI1_RXPOLARITY_0_net), 
        .RXSTANDBYSTATUS_0(
        PCIE_1_RXSTANDBYSTATUS_2_PCIESS_LANE2_Pipe_AXI1_RXSTANDBYSTATUS_0_net)
        , .RXSTATUS_0({
        PCIE_1_RXSTATUS_2_PCIESS_LANE2_Pipe_AXI1_RXSTATUS_0_net_2, 
        PCIE_1_RXSTATUS_2_PCIESS_LANE2_Pipe_AXI1_RXSTATUS_0_net_1, 
        PCIE_1_RXSTATUS_2_PCIESS_LANE2_Pipe_AXI1_RXSTATUS_0_net_0}), 
        .RXVALID_0(
        PCIE_1_RXVALID_2_PCIESS_LANE2_Pipe_AXI1_RXVALID_0_net), 
        .TXCOMPLIANCE_0(
        PCIE_1_TXCOMPLIANCE_2_PCIESS_LANE2_Pipe_AXI1_TXCOMPLIANCE_0_net)
        , .TXDATA_0({
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_31, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_30, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_29, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_28, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_27, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_26, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_25, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_24, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_23, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_22, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_21, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_20, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_19, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_18, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_17, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_16, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_15, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_14, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_13, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_12, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_11, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_10, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_9, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_8, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_7, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_6, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_5, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_4, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_3, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_2, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_1, 
        PCIE_1_TXDATA_2_PCIESS_LANE2_Pipe_AXI1_TXDATA_0_net_0}), 
        .TXDATAK_0({
        PCIE_1_TXDATAK_2_PCIESS_LANE2_Pipe_AXI1_TXDATAK_0_net_3, 
        PCIE_1_TXDATAK_2_PCIESS_LANE2_Pipe_AXI1_TXDATAK_0_net_2, 
        PCIE_1_TXDATAK_2_PCIESS_LANE2_Pipe_AXI1_TXDATAK_0_net_1, 
        PCIE_1_TXDATAK_2_PCIESS_LANE2_Pipe_AXI1_TXDATAK_0_net_0}), 
        .TXDATAVALID_0(
        PCIE_1_TXDATAVALID_2_PCIESS_LANE2_Pipe_AXI1_TXDATAVALID_0_net), 
        .TXDEEMPH(PCIE_1_TXDEEMPH_PCIESS_LANE2_Pipe_AXI1_TXDEEMPH_net), 
        .TXDETECTRX_LOOPBACK_0(
        PCIE_1_TXDETECTRX_LOOPBACK_2_PCIESS_LANE2_Pipe_AXI1_TXDETECTRX_LOOPBACK_0_net)
        , .TXELECIDLE_0(
        PCIE_1_TXELECIDLE_2_PCIESS_LANE2_Pipe_AXI1_TXELECIDLE_0_net), 
        .TXMARGIN({
        PCIE_1_TXMARGIN_PCIESS_LANE2_Pipe_AXI1_TXMARGIN_net_2, 
        PCIE_1_TXMARGIN_PCIESS_LANE2_Pipe_AXI1_TXMARGIN_net_1, 
        PCIE_1_TXMARGIN_PCIESS_LANE2_Pipe_AXI1_TXMARGIN_net_0}), 
        .TXSWING(PCIE_1_TXSWING_PCIESS_LANE2_Pipe_AXI1_TXSWING_net), 
        .PIPE_CLK_0(
        PCIE_1_PIPE_CLK_2_PCIESS_LANE2_Pipe_AXI1_PIPE_CLK_0_net), 
        .PCLK_OUT_0(
        PCIE_1_PCLK_OUT_2_PCIESS_LANE2_Pipe_AXI1_PCLK_OUT_0_net), 
        .AXI_CLK(PCIE_COMMON_AXI_CLK_OUT_net), .LINK_CLK(gnd_net), 
        .LINK_ADDR({gnd_net, gnd_net, gnd_net}), .LINK_EN(gnd_net), 
        .LINK_ARST_N(gnd_net), .LINK_WDATA({gnd_net, gnd_net, gnd_net, 
        gnd_net}), .LINK_RDATA({nc380, nc381, nc382, nc383}));
    GND PCIESS_AXI_1_M_AWID_3_GndInst (.Y(PCIESS_AXI_1_M_AWID[3]));
    XCVR_APB_LINK pcie_apblink_inst (.S_RDATA({
        pcie_apblink_master_inst_lnk_m_rdata_pcie_apblink_inst_S_RDATA_net_3, 
        pcie_apblink_master_inst_lnk_m_rdata_pcie_apblink_inst_S_RDATA_net_2, 
        pcie_apblink_master_inst_lnk_m_rdata_pcie_apblink_inst_S_RDATA_net_1, 
        pcie_apblink_master_inst_lnk_m_rdata_pcie_apblink_inst_S_RDATA_net_0})
        , .S_ADDR({
        pcie_apblink_master_inst_lnk_m_addr_pcie_apblink_inst_S_ADDR_net_2, 
        pcie_apblink_master_inst_lnk_m_addr_pcie_apblink_inst_S_ADDR_net_1, 
        pcie_apblink_master_inst_lnk_m_addr_pcie_apblink_inst_S_ADDR_net_0})
        , .S_CLK(
        pcie_apblink_master_inst_lnk_m_clock_pcie_apblink_inst_S_CLK_net)
        , .S_EN(
        pcie_apblink_master_inst_lnk_m_enable_pcie_apblink_inst_S_EN_net)
        , .S_ARST_N(
        pcie_apblink_master_inst_lnk_m_rst_b_pcie_apblink_inst_S_ARST_N_net)
        , .S_WDATA({
        pcie_apblink_master_inst_lnk_m_wdata_pcie_apblink_inst_S_WDATA_net_3, 
        pcie_apblink_master_inst_lnk_m_wdata_pcie_apblink_inst_S_WDATA_net_2, 
        pcie_apblink_master_inst_lnk_m_wdata_pcie_apblink_inst_S_WDATA_net_1, 
        pcie_apblink_master_inst_lnk_m_wdata_pcie_apblink_inst_S_WDATA_net_0})
        , .PCIE0_BRIDGE_CLK(), .PCIE0_BRIDGE_ADDR({nc384, nc385, nc386})
        , .PCIE0_BRIDGE_EN(), .PCIE0_BRIDGE_ARST_N(), 
        .PCIE0_BRIDGE_WDATA({nc387, nc388, nc389, nc390}), 
        .PCIE0_BRIDGE_RDATA({nc391, nc392, nc393, nc394}), 
        .PCIE0_CTRL_CLK(), .PCIE0_CTRL_ADDR({nc395, nc396, nc397}), 
        .PCIE0_CTRL_EN(), .PCIE0_CTRL_ARST_N(), .PCIE0_CTRL_WDATA({
        nc398, nc399, nc400, nc401}), .PCIE0_CTRL_RDATA({nc402, nc403, 
        nc404, nc405}), .PCIE1_BRIDGE_CLK(
        pcie_apblink_inst_PCIE1_BRIDGE_CLK_PCIE_1_LINK_BRIDGE_CLK_net), 
        .PCIE1_BRIDGE_ADDR({
        pcie_apblink_inst_PCIE1_BRIDGE_ADDR_PCIE_1_LINK_BRIDGE_ADDR_net_2, 
        pcie_apblink_inst_PCIE1_BRIDGE_ADDR_PCIE_1_LINK_BRIDGE_ADDR_net_1, 
        pcie_apblink_inst_PCIE1_BRIDGE_ADDR_PCIE_1_LINK_BRIDGE_ADDR_net_0})
        , .PCIE1_BRIDGE_EN(
        pcie_apblink_inst_PCIE1_BRIDGE_EN_PCIE_1_LINK_BRIDGE_EN_net), 
        .PCIE1_BRIDGE_ARST_N(
        pcie_apblink_inst_PCIE1_BRIDGE_ARST_N_PCIE_1_LINK_BRIDGE_ARST_N_net)
        , .PCIE1_BRIDGE_WDATA({
        pcie_apblink_inst_PCIE1_BRIDGE_WDATA_PCIE_1_LINK_BRIDGE_WDATA_net_3, 
        pcie_apblink_inst_PCIE1_BRIDGE_WDATA_PCIE_1_LINK_BRIDGE_WDATA_net_2, 
        pcie_apblink_inst_PCIE1_BRIDGE_WDATA_PCIE_1_LINK_BRIDGE_WDATA_net_1, 
        pcie_apblink_inst_PCIE1_BRIDGE_WDATA_PCIE_1_LINK_BRIDGE_WDATA_net_0})
        , .PCIE1_BRIDGE_RDATA({
        pcie_apblink_inst_PCIE1_BRIDGE_RDATA_PCIE_1_LINK_BRIDGE_RDATA_net_3, 
        pcie_apblink_inst_PCIE1_BRIDGE_RDATA_PCIE_1_LINK_BRIDGE_RDATA_net_2, 
        pcie_apblink_inst_PCIE1_BRIDGE_RDATA_PCIE_1_LINK_BRIDGE_RDATA_net_1, 
        pcie_apblink_inst_PCIE1_BRIDGE_RDATA_PCIE_1_LINK_BRIDGE_RDATA_net_0})
        , .PCIE1_CTRL_CLK(), .PCIE1_CTRL_ADDR({nc406, nc407, nc408}), 
        .PCIE1_CTRL_EN(), .PCIE1_CTRL_ARST_N(), .PCIE1_CTRL_WDATA({
        nc409, nc410, nc411, nc412}), .PCIE1_CTRL_RDATA({nc413, nc414, 
        nc415, nc416}), .EXT_PLL_0_CLK(), .EXT_PLL_0_ADDR({nc417, 
        nc418, nc419}), .EXT_PLL_0_EN(), .EXT_PLL_0_ARST_N(), 
        .EXT_PLL_0_WDATA({nc420, nc421, nc422, nc423}), 
        .EXT_PLL_0_RDATA({gnd_net, gnd_net, gnd_net, gnd_net}), 
        .EXT_PLL_1_CLK(), .EXT_PLL_1_ADDR({nc424, nc425, nc426}), 
        .EXT_PLL_1_EN(), .EXT_PLL_1_ARST_N(), .EXT_PLL_1_WDATA({nc427, 
        nc428, nc429, nc430}), .EXT_PLL_1_RDATA({gnd_net, gnd_net, 
        gnd_net, gnd_net}), .QUAD_PLL_CLK(), .QUAD_PLL_ADDR({nc431, 
        nc432, nc433}), .QUAD_PLL_EN(), .QUAD_PLL_ARST_N(), 
        .QUAD_PLL_WDATA({nc434, nc435, nc436, nc437}), .QUAD_PLL_RDATA({
        gnd_net, gnd_net, gnd_net, gnd_net}), .L0_CLK(), .L0_ADDR({
        nc438, nc439, nc440}), .L0_EN(), .L0_ARST_N(), .L0_WDATA({
        nc441, nc442, nc443, nc444}), .L0_RDATA({gnd_net, gnd_net, 
        gnd_net, gnd_net}), .L1_CLK(), .L1_ADDR({nc445, nc446, nc447}), 
        .L1_EN(), .L1_ARST_N(), .L1_WDATA({nc448, nc449, nc450, nc451})
        , .L1_RDATA({gnd_net, gnd_net, gnd_net, gnd_net}), .L2_CLK(), 
        .L2_ADDR({nc452, nc453, nc454}), .L2_EN(), .L2_ARST_N(), 
        .L2_WDATA({nc455, nc456, nc457, nc458}), .L2_RDATA({gnd_net, 
        gnd_net, gnd_net, gnd_net}), .L3_CLK(), .L3_ADDR({nc459, nc460, 
        nc461}), .L3_EN(), .L3_ARST_N(), .L3_WDATA({nc462, nc463, 
        nc464, nc465}), .L3_RDATA({gnd_net, gnd_net, gnd_net, gnd_net})
        );
    GND PCIESS_AXI_1_M_ARLEN_7_GndInst (.Y(PCIESS_AXI_1_M_ARLEN[7]));
    
endmodule
